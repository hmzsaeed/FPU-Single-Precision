##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Tue May 31 01:06:29 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_proj_example
  CLASS BLOCK ;
  SIZE 929.200000 BY 920.720000 ;
  FOREIGN user_proj_example 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.852 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.613 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 131.062 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 699.936 LAYER met3  ;
    ANTENNAGATEAREA 0.852 LAYER met3  ;
    ANTENNAMAXAREACAR 154.522 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 823.871 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.107277 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1.830000 0.000000 1.970000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2375 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.161 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.1466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 263.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2275 LAYER met4  ;
    ANTENNAMAXAREACAR 24.4366 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 126.994 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.243591 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 4.180000 0.490000 4.320000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.530000 0.000000 197.670000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.430000 0.000000 66.570000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.430000 0.000000 199.570000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.630000 0.000000 195.770000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.730000 0.000000 193.870000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.830000 0.000000 191.970000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.930000 0.000000 190.070000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.230000 0.000000 127.370000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.330000 0.000000 125.470000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.430000 0.000000 123.570000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530000 0.000000 121.670000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.630000 0.000000 119.770000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.730000 0.000000 117.870000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.830000 0.000000 115.970000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.930000 0.000000 114.070000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.030000 0.000000 112.170000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.130000 0.000000 110.270000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.230000 0.000000 108.370000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.330000 0.000000 106.470000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.430000 0.000000 104.570000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.530000 0.000000 102.670000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.630000 0.000000 100.770000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.730000 0.000000 98.870000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.830000 0.000000 96.970000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.930000 0.000000 95.070000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.030000 0.000000 93.170000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.130000 0.000000 91.270000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.230000 0.000000 89.370000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.330000 0.000000 87.470000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.430000 0.000000 85.570000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.530000 0.000000 83.670000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.630000 0.000000 81.770000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.730000 0.000000 79.870000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830000 0.000000 77.970000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.930000 0.000000 76.070000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.030000 0.000000 74.170000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.130000 0.000000 72.270000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.230000 0.000000 70.370000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.330000 0.000000 68.470000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.530000 0.000000 64.670000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.630000 0.000000 62.770000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.730000 0.000000 60.870000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.830000 0.000000 58.970000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.930000 0.000000 57.070000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.030000 0.000000 55.170000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.130000 0.000000 53.270000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.230000 0.000000 51.370000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.330000 0.000000 49.470000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.430000 0.000000 47.570000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.530000 0.000000 45.670000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.630000 0.000000 43.770000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.730000 0.000000 41.870000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.830000 0.000000 39.970000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.930000 0.000000 38.070000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.030000 0.000000 36.170000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130000 0.000000 34.270000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.230000 0.000000 32.370000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.330000 0.000000 30.470000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.430000 0.000000 28.570000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.530000 0.000000 26.670000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.630000 0.000000 24.770000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.730000 0.000000 22.870000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.830000 0.000000 20.970000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.930000 0.000000 19.070000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.030000 0.000000 17.170000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.130000 0.000000 15.270000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.230000 0.000000 13.370000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.330000 0.000000 11.470000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.430000 0.000000 9.570000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.530000 0.000000 7.670000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.630000 0.000000 5.770000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 3.730000 0.000000 3.870000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 188.030000 0.000000 188.170000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 186.130000 0.000000 186.270000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.714 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 184.230000 0.000000 184.370000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 182.330000 0.000000 182.470000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 180.430000 0.000000 180.570000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.714 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 178.530000 0.000000 178.670000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.714 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 176.630000 0.000000 176.770000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.714 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 174.730000 0.000000 174.870000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.714 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 172.830000 0.000000 172.970000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 170.930000 0.000000 171.070000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 169.030000 0.000000 169.170000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 167.130000 0.000000 167.270000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 165.230000 0.000000 165.370000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 163.330000 0.000000 163.470000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 161.430000 0.000000 161.570000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 159.530000 0.000000 159.670000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 157.630000 0.000000 157.770000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 155.730000 0.000000 155.870000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 153.830000 0.000000 153.970000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 151.930000 0.000000 152.070000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 150.030000 0.000000 150.170000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 148.130000 0.000000 148.270000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 146.230000 0.000000 146.370000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 144.330000 0.000000 144.470000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 142.430000 0.000000 142.570000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 140.530000 0.000000 140.670000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 138.630000 0.000000 138.770000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 136.730000 0.000000 136.870000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.714 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 134.830000 0.000000 134.970000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.714 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 132.930000 0.000000 133.070000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 131.030000 0.000000 131.170000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3358 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.518 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 129.130000 0.000000 129.270000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.630000 0.000000 442.770000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.730000 0.000000 440.870000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.830000 0.000000 438.970000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.930000 0.000000 437.070000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.030000 0.000000 435.170000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.130000 0.000000 433.270000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.230000 0.000000 431.370000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.330000 0.000000 429.470000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430000 0.000000 427.570000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.530000 0.000000 425.670000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.630000 0.000000 423.770000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.730000 0.000000 421.870000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.830000 0.000000 419.970000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.930000 0.000000 418.070000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.030000 0.000000 416.170000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.130000 0.000000 414.270000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.230000 0.000000 412.370000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.330000 0.000000 410.470000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.430000 0.000000 408.570000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.530000 0.000000 406.670000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.630000 0.000000 404.770000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.730000 0.000000 402.870000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.830000 0.000000 400.970000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.930000 0.000000 399.070000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.030000 0.000000 397.170000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.130000 0.000000 395.270000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.230000 0.000000 393.370000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.330000 0.000000 391.470000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.430000 0.000000 389.570000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.530000 0.000000 387.670000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.630000 0.000000 385.770000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730000 0.000000 383.870000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.830000 0.000000 381.970000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.930000 0.000000 380.070000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.030000 0.000000 378.170000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.130000 0.000000 376.270000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.230000 0.000000 374.370000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.330000 0.000000 372.470000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.430000 0.000000 370.570000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.530000 0.000000 368.670000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.630000 0.000000 366.770000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730000 0.000000 364.870000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.830000 0.000000 362.970000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.930000 0.000000 361.070000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.030000 0.000000 359.170000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.130000 0.000000 357.270000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.230000 0.000000 355.370000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.330000 0.000000 353.470000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.430000 0.000000 351.570000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.530000 0.000000 349.670000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.630000 0.000000 347.770000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.730000 0.000000 345.870000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.830000 0.000000 343.970000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.930000 0.000000 342.070000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030000 0.000000 340.170000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.130000 0.000000 338.270000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.230000 0.000000 336.370000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.330000 0.000000 334.470000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.430000 0.000000 332.570000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.530000 0.000000 330.670000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.630000 0.000000 328.770000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.730000 0.000000 326.870000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.434 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 68.3778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 365.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.94 LAYER met4  ;
    ANTENNAMAXAREACAR 14.617 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 73.9351 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.221145 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 324.830000 0.000000 324.970000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3583 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 255.835 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1370.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 14.9265 LAYER met4  ;
    ANTENNAMAXAREACAR 65.9874 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 333.061 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 322.930000 0.000000 323.070000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.030000 0.000000 321.170000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.130000 0.000000 319.270000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.230000 0.000000 317.370000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.330000 0.000000 315.470000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.430000 0.000000 313.570000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.530000 0.000000 311.670000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.630000 0.000000 309.770000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.730000 0.000000 307.870000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.830000 0.000000 305.970000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.930000 0.000000 304.070000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.030000 0.000000 302.170000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.130000 0.000000 300.270000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.230000 0.000000 298.370000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330000 0.000000 296.470000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.430000 0.000000 294.570000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.530000 0.000000 292.670000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.630000 0.000000 290.770000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.730000 0.000000 288.870000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.830000 0.000000 286.970000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.930000 0.000000 285.070000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.030000 0.000000 283.170000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.130000 0.000000 281.270000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.230000 0.000000 279.370000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.330000 0.000000 277.470000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.430000 0.000000 275.570000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.530000 0.000000 273.670000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.630000 0.000000 271.770000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.730000 0.000000 269.870000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.830000 0.000000 267.970000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.930000 0.000000 266.070000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.030000 0.000000 264.170000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.130000 0.000000 262.270000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.493 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 18.5058 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 87.7309 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.137617 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 260.230000 0.000000 260.370000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.47 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.124 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met2  ;
    ANTENNAMAXAREACAR 3.9371 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.6498 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0735354 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 258.330000 0.000000 258.470000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0486 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.017 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 14.053 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.8727 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 256.430000 0.000000 256.570000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.544 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2275 LAYER met2  ;
    ANTENNAMAXAREACAR 2.33001 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.90617 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 254.530000 0.000000 254.670000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0912 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.122 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 6.03212 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.3313 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 252.630000 0.000000 252.770000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7488 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.636 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 6.73992 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.1507 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.134949 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 250.730000 0.000000 250.870000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.4328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.112 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 24.6304 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 126.421 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 248.830000 0.000000 248.970000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7376 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.354 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 5.83907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.2921 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 246.930000 0.000000 247.070000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.514 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 20.5309 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 99.7232 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 245.030000 0.000000 245.170000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4084 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.816 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 19.0989 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 91.716 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 243.130000 0.000000 243.270000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.12 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.567 LAYER met2  ;
    ANTENNAMAXAREACAR 7.12555 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.4782 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.203968 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 241.230000 0.000000 241.370000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.71 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2275 LAYER met2  ;
    ANTENNAMAXAREACAR 3.60314 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.4334 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.330000 0.000000 239.470000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.5908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met3  ;
    ANTENNAMAXAREACAR 11.8937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 61.3665 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.24 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 237.430000 0.000000 237.570000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.969 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 8.44903 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.8222 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 235.530000 0.000000 235.670000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6667 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.0528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met3  ;
    ANTENNAMAXAREACAR 7.57366 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 32.7838 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.24 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 233.630000 0.000000 233.770000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met2  ;
    ANTENNAMAXAREACAR 5.05091 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.2761 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.162222 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 231.730000 0.000000 231.870000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.830000 0.000000 229.970000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.930000 0.000000 228.070000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.030000 0.000000 226.170000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.130000 0.000000 224.270000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.230000 0.000000 222.370000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.330000 0.000000 220.470000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.430000 0.000000 218.570000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.530000 0.000000 216.670000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.630000 0.000000 214.770000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.730000 0.000000 212.870000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.830000 0.000000 210.970000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930000 0.000000 209.070000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.030000 0.000000 207.170000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.130000 0.000000 205.270000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.053 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.803 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 20.2359 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.9293 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 203.230000 0.000000 203.370000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.330000 0.000000 201.470000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.342 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 685.830000 0.000000 685.970000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 683.930000 0.000000 684.070000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 682.030000 0.000000 682.170000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 680.130000 0.000000 680.270000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 678.230000 0.000000 678.370000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 676.330000 0.000000 676.470000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 674.430000 0.000000 674.570000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 672.530000 0.000000 672.670000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 670.630000 0.000000 670.770000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 668.730000 0.000000 668.870000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 666.830000 0.000000 666.970000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 664.930000 0.000000 665.070000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 663.030000 0.000000 663.170000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 661.130000 0.000000 661.270000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 659.230000 0.000000 659.370000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 657.330000 0.000000 657.470000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 655.430000 0.000000 655.570000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 653.530000 0.000000 653.670000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 651.630000 0.000000 651.770000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 649.730000 0.000000 649.870000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 647.830000 0.000000 647.970000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 645.930000 0.000000 646.070000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 644.030000 0.000000 644.170000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 642.130000 0.000000 642.270000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 640.230000 0.000000 640.370000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 638.330000 0.000000 638.470000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 636.430000 0.000000 636.570000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 634.530000 0.000000 634.670000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 632.630000 0.000000 632.770000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 630.730000 0.000000 630.870000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 628.830000 0.000000 628.970000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 626.930000 0.000000 627.070000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 625.030000 0.000000 625.170000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 623.130000 0.000000 623.270000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 621.230000 0.000000 621.370000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 619.330000 0.000000 619.470000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 617.430000 0.000000 617.570000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 615.530000 0.000000 615.670000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 613.630000 0.000000 613.770000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 611.730000 0.000000 611.870000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 609.830000 0.000000 609.970000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 607.930000 0.000000 608.070000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 606.030000 0.000000 606.170000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 604.130000 0.000000 604.270000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 602.230000 0.000000 602.370000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 600.330000 0.000000 600.470000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 598.430000 0.000000 598.570000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 596.530000 0.000000 596.670000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 594.630000 0.000000 594.770000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 592.730000 0.000000 592.870000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 590.830000 0.000000 590.970000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 588.930000 0.000000 589.070000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 587.030000 0.000000 587.170000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 585.130000 0.000000 585.270000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 583.230000 0.000000 583.370000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 581.330000 0.000000 581.470000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 579.430000 0.000000 579.570000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 577.530000 0.000000 577.670000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 575.630000 0.000000 575.770000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 573.730000 0.000000 573.870000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 571.830000 0.000000 571.970000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 569.930000 0.000000 570.070000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 568.030000 0.000000 568.170000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.342 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 566.130000 0.000000 566.270000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.574 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.439 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 96.3768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 514.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 564.230000 0.000000 564.370000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 89.9718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 480.32 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 562.330000 0.000000 562.470000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7185 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 92.3508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 493.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 560.430000 0.000000 560.570000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.6908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 473.488 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 558.530000 0.000000 558.670000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.7038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 484.224 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 556.630000 0.000000 556.770000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8181 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 92.7168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 494.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 554.730000 0.000000 554.870000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 92.8998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 495.936 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 552.830000 0.000000 552.970000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8211 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 97.8408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 522.288 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 550.930000 0.000000 551.070000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.0025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.1418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 470.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 549.030000 0.000000 549.170000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5274 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.476 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.4436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 472.64 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 547.130000 0.000000 547.270000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 93.4488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 498.864 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 545.230000 0.000000 545.370000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8543 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 87.7998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 468.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 543.330000 0.000000 543.470000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7357 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.3378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 482.272 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 541.430000 0.000000 541.570000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5757 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.4436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 472.64 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 539.530000 0.000000 539.670000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3415 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.3248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 471.536 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 537.630000 0.000000 537.770000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 82.8348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 442.256 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 535.730000 0.000000 535.870000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7469 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 96.5598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 515.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 533.830000 0.000000 533.970000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 87.0438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 464.704 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 531.930000 0.000000 532.070000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 86.8608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 463.728 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 530.030000 0.000000 530.170000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5865 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.403 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 89.7888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 479.344 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 528.130000 0.000000 528.270000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7141 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.4095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.713 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5445 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.1418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 470.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 526.230000 0.000000 526.370000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6639 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.6908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 473.488 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 524.330000 0.000000 524.470000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.6565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 84.6648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 452.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 522.430000 0.000000 522.570000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8515 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 87.4098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 466.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 520.530000 0.000000 520.670000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4073 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.0776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 470.688 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 518.630000 0.000000 518.770000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 86.9634 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 465.216 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 516.730000 0.000000 516.870000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 91.0698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 486.176 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 514.830000 0.000000 514.970000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7749 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 89.2302 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 477.776 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 512.930000 0.000000 513.070000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5977 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.412 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 85.7628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 457.872 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 511.030000 0.000000 511.170000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.8745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 74.3526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 397.488 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 509.130000 0.000000 509.270000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7357 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 85.5798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 456.896 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 507.230000 0.000000 507.370000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2409 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 91.8018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 490.08 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 505.330000 0.000000 505.470000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.492 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 503.430000 0.000000 503.570000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 501.530000 0.000000 501.670000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 499.630000 0.000000 499.770000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 497.730000 0.000000 497.870000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 495.830000 0.000000 495.970000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 493.930000 0.000000 494.070000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 492.030000 0.000000 492.170000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 490.130000 0.000000 490.270000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 488.230000 0.000000 488.370000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 486.330000 0.000000 486.470000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 484.430000 0.000000 484.570000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 482.530000 0.000000 482.670000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 480.630000 0.000000 480.770000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 478.730000 0.000000 478.870000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 476.830000 0.000000 476.970000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 474.930000 0.000000 475.070000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 473.030000 0.000000 473.170000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 471.130000 0.000000 471.270000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 469.230000 0.000000 469.370000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 467.330000 0.000000 467.470000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 465.430000 0.000000 465.570000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 463.530000 0.000000 463.670000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 461.630000 0.000000 461.770000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 459.730000 0.000000 459.870000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.443 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 457.830000 0.000000 457.970000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 455.930000 0.000000 456.070000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 454.030000 0.000000 454.170000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 452.130000 0.000000 452.270000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 450.230000 0.000000 450.370000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 448.330000 0.000000 448.470000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 446.430000 0.000000 446.570000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 444.530000 0.000000 444.670000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.030000 0.000000 929.170000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.130000 0.000000 927.270000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.230000 0.000000 925.370000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.330000 0.000000 923.470000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.430000 0.000000 921.570000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.530000 0.000000 919.670000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.630000 0.000000 917.770000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.730000 0.000000 915.870000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.830000 0.000000 913.970000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.930000 0.000000 912.070000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.030000 0.000000 910.170000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130000 0.000000 908.270000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.230000 0.000000 906.370000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.330000 0.000000 904.470000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.430000 0.000000 902.570000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.530000 0.000000 900.670000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.630000 0.000000 898.770000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.730000 0.000000 896.870000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.830000 0.000000 894.970000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.930000 0.000000 893.070000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.030000 0.000000 891.170000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130000 0.000000 889.270000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.230000 0.000000 887.370000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.330000 0.000000 885.470000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.430000 0.000000 883.570000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.530000 0.000000 881.670000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.630000 0.000000 879.770000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.730000 0.000000 877.870000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.830000 0.000000 875.970000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.930000 0.000000 874.070000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.030000 0.000000 872.170000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.130000 0.000000 870.270000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.230000 0.000000 868.370000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.330000 0.000000 866.470000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.430000 0.000000 864.570000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.530000 0.000000 862.670000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.630000 0.000000 860.770000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.730000 0.000000 858.870000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.830000 0.000000 856.970000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.930000 0.000000 855.070000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.030000 0.000000 853.170000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.130000 0.000000 851.270000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.230000 0.000000 849.370000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.330000 0.000000 847.470000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.430000 0.000000 845.570000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.530000 0.000000 843.670000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.630000 0.000000 841.770000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.730000 0.000000 839.870000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.830000 0.000000 837.970000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.930000 0.000000 836.070000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.030000 0.000000 834.170000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.130000 0.000000 832.270000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.230000 0.000000 830.370000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.330000 0.000000 828.470000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.430000 0.000000 826.570000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.530000 0.000000 824.670000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.630000 0.000000 822.770000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730000 0.000000 820.870000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.830000 0.000000 818.970000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.930000 0.000000 817.070000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.030000 0.000000 815.170000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.130000 0.000000 813.270000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5573 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 72.7698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 388.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.94 LAYER met4  ;
    ANTENNAMAXAREACAR 14.0324 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 72.7481 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0832155 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 811.230000 0.000000 811.370000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.9389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 144.189 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2185 LAYER met2  ;
    ANTENNAMAXAREACAR 19.0358 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 91.2281 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.0875366 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 2.2185 LAYER met3  ;
    ANTENNAMAXAREACAR 19.1489 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 92.043 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.105567 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 199.82 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1068.99 LAYER met4  ;
    ANTENNAGATEAREA 22.7625 LAYER met4  ;
    ANTENNAMAXAREACAR 59.1856 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 301.399 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521429 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 809.330000 0.000000 809.470000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.91 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.1175 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.0992 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 807.430000 0.000000 807.570000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.323 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.9361 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.8929 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 805.530000 0.000000 805.670000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.169 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 16.4135 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.5992 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 803.630000 0.000000 803.770000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7114 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.449 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.1222 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.3452 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 801.730000 0.000000 801.870000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6344 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.3397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.2103 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 799.830000 0.000000 799.970000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.1583 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.004 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 797.930000 0.000000 798.070000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.337 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.0762 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.377 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 796.030000 0.000000 796.170000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9095 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 21.5167 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.3175 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 794.130000 0.000000 794.270000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6008 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.896 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.0952 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.9881 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 792.230000 0.000000 792.370000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.547 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.2917 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.6706 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 790.330000 0.000000 790.470000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.183 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 16.4357 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.7103 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 788.430000 0.000000 788.570000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7142 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.463 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.1444 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.4564 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 786.530000 0.000000 786.670000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.707 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 16.773 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.377 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 784.630000 0.000000 784.770000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.141 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 16.7401 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.4484 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 782.730000 0.000000 782.870000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7394 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.589 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.9873 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.9325 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 780.830000 0.000000 780.970000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6358 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.071 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 19.0556 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.0119 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 778.930000 0.000000 779.070000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.861 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 16.1103 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.5992 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 777.030000 0.000000 777.170000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.717 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.477 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.2734 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.1151 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 775.130000 0.000000 775.270000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7086 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.435 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.7651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.8214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 773.230000 0.000000 773.370000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.239 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 19.8333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.9008 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 771.330000 0.000000 771.470000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5826 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.805 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 16.9286 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.1548 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 769.430000 0.000000 769.570000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.799 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 19.7139 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.7817 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 767.530000 0.000000 767.670000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7422 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.603 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 20.5651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 91.8214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 765.630000 0.000000 765.770000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.4988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.464 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 16.4722 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 79.6032 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 763.730000 0.000000 763.870000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.847 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.5063 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.0436 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 761.830000 0.000000 761.970000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.169 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.6917 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.6706 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 759.930000 0.000000 760.070000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7114 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.449 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 20.3206 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.5992 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 758.030000 0.000000 758.170000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.577 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.777 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 22.4444 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 101.956 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 756.130000 0.000000 756.270000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.679 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.2619 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.8214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 754.230000 0.000000 754.370000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.337 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.0512 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.004 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 752.330000 0.000000 752.470000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.745 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.617 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 19.5651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.8214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 750.430000 0.000000 750.570000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.575 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 22.4111 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 101.79 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 748.530000 0.000000 748.670000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7142 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.463 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met2  ;
    ANTENNAMAXAREACAR 2.02628 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.2895 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0446181 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 746.630000 0.000000 746.770000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9914 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.849 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met2  ;
    ANTENNAMAXAREACAR 2.58974 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.0482 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0446181 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 744.730000 0.000000 744.870000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6666 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.225 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met2  ;
    ANTENNAMAXAREACAR 1.98496 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.0829 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0446181 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 742.830000 0.000000 742.970000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.121 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.304 LAYER met2  ;
    ANTENNAMAXAREACAR 1.94967 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.66168 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.022309 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 740.930000 0.000000 741.070000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0166 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.975 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met2  ;
    ANTENNAMAXAREACAR 2.28878 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.602 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0446181 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 739.030000 0.000000 739.170000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.351 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.576 LAYER met2  ;
    ANTENNAMAXAREACAR 3.625 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.0391 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0892361 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 737.130000 0.000000 737.270000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6974 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.379 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 3.84162 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.3707 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 735.230000 0.000000 735.370000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4058 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.921 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met2  ;
    ANTENNAMAXAREACAR 2.62663 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.2912 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0446181 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 733.330000 0.000000 733.470000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.576 LAYER met2  ;
    ANTENNAMAXAREACAR 3.75538 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.5738 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0892361 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 731.430000 0.000000 731.570000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.661 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.197 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 3.76808 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.003 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 729.530000 0.000000 729.670000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6638 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.211 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met2  ;
    ANTENNAMAXAREACAR 1.98253 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.07075 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0446181 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 727.630000 0.000000 727.770000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.947 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met2  ;
    ANTENNAMAXAREACAR 2.28392 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.57769 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0446181 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 725.730000 0.000000 725.870000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.127 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 3.7398 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.8616 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 723.830000 0.000000 723.970000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.085 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 3.82364 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.1444 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 721.930000 0.000000 722.070000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6344 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.576 LAYER met2  ;
    ANTENNAMAXAREACAR 3.71649 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.3793 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0892361 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 720.030000 0.000000 720.170000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7418 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.601 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met2  ;
    ANTENNAMAXAREACAR 3.07342 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.4666 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0446181 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 718.130000 0.000000 718.270000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.230000 0.000000 716.370000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.330000 0.000000 714.470000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.430000 0.000000 712.570000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.530000 0.000000 710.670000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.630000 0.000000 708.770000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.730000 0.000000 706.870000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.830000 0.000000 704.970000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.930000 0.000000 703.070000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.030000 0.000000 701.170000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.130000 0.000000 699.270000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.230000 0.000000 697.370000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.330000 0.000000 695.470000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.430000 0.000000 693.570000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.530000 0.000000 691.670000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 8.43333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.3646 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 689.630000 0.000000 689.770000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.730000 0.000000 687.870000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 44.760000 0.800000 45.060000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 112.130000 0.800000 112.430000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 179.500000 0.800000 179.800000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 246.865000 0.800000 247.165000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 314.235000 0.800000 314.535000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 381.600000 0.800000 381.900000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 448.970000 0.800000 449.270000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 516.340000 0.800000 516.640000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 583.705000 0.800000 584.005000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 651.075000 0.800000 651.375000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 718.440000 0.800000 718.740000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 785.810000 0.800000 786.110000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 853.180000 0.800000 853.480000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 913.020000 0.800000 913.320000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.405000 920.230000 71.545000 920.720000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.620000 920.230000 178.760000 920.720000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.835000 920.230000 285.975000 920.720000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.050000 920.230000 393.190000 920.720000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.260000 920.230000 500.400000 920.720000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.475000 920.230000 607.615000 920.720000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.690000 920.230000 714.830000 920.720000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.905000 920.230000 822.045000 920.720000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.560000 920.230000 915.700000 920.720000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 878.700000 929.200000 879.000000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 815.925000 929.200000 816.225000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 753.150000 929.200000 753.450000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 690.375000 929.200000 690.675000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 627.600000 929.200000 627.900000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 564.825000 929.200000 565.125000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 502.050000 929.200000 502.350000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 439.275000 929.200000 439.575000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 376.500000 929.200000 376.800000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2979 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 13.8756 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 64.9414 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 313.725000 929.200000 314.025000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 250.950000 929.200000 251.250000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 188.175000 929.200000 188.475000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 125.400000 929.200000 125.700000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 62.625000 929.200000 62.925000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.400000 9.610000 929.200000 9.910000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.353 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.99 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.519 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 22.305000 0.800000 22.605000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 99.7561 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 532.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 65.0196 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 347.712 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 89.675000 0.800000 89.975000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.5374 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 173.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.8026 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.888 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 157.040000 0.800000 157.340000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 117.941 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 629.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.3468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.32 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 224.410000 0.800000 224.710000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 156.544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 835.368 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 291.780000 0.800000 292.080000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 136.544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 728.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.1508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.608 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 359.145000 0.800000 359.445000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 154.66 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 825.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.2558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.168 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 426.515000 0.800000 426.815000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 151.068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 806.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.8308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 63.568 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 493.880000 0.800000 494.180000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 139.557 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 744.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.2748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.936 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 561.250000 0.800000 561.550000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 128.271 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 684.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.1056 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 193.504 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 628.620000 0.800000 628.920000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 83.7199 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 446.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.8966 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 171.056 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 695.985000 0.800000 696.285000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 147.692 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 788.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.9478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 160.192 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 763.355000 0.800000 763.655000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 118.974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 634.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.0328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.312 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 830.720000 0.800000 831.020000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 63.8251 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 341.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.8056 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.904 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 898.090000 0.800000 898.390000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.0457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.0675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 60.0658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 321.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.5964 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 276.592 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 35.670000 920.230000 35.810000 920.720000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6019 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.8485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.978 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 283.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 138.101 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 737.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 142.880000 920.230000 143.020000 920.720000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4853 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.2655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 147.553 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 787.888 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 250.095000 920.230000 250.235000 920.720000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.9771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.7245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 125.474 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 669.664 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 357.310000 920.230000 357.450000 920.720000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.6028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.5106 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 227.664 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 464.525000 920.230000 464.665000 920.720000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.7138 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 132.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.0978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 208.992 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 571.740000 920.230000 571.880000 920.720000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.6371 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 147.906 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 74.0508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 395.408 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 678.950000 920.230000 679.090000 920.720000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3676 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.526 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 84.2128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 450.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.0068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 786.165000 920.230000 786.305000 920.720000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1655 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 90.5368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 483.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.4118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 168 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 893.380000 920.230000 893.520000 920.720000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 93.2449 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.2478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 257.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 899.625000 929.200000 899.925000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.1194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.9408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.488 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 836.850000 929.200000 837.150000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 93.3499 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 498.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.8298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 212.896 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 774.075000 929.200000 774.375000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 122.57 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 655.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 112.607 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 601.984 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 711.300000 929.200000 711.600000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 113.862 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 608.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.7918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.36 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 648.525000 929.200000 648.825000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 123.193 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 657.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 69.2526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 370.288 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 585.750000 929.200000 586.050000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.2284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 114.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.9418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.16 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 522.975000 929.200000 523.275000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 118.821 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 634.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.2298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.696 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 460.200000 929.200000 460.500000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3991 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.4466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.656 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 397.425000 929.200000 397.725000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.37 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.68 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.531 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 334.650000 929.200000 334.950000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7101 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.9834 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.656 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 271.875000 929.200000 272.175000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 209.100000 929.200000 209.400000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 146.325000 929.200000 146.625000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.37 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.68 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.531 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 83.550000 929.200000 83.850000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.37 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.68 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.531 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 20.775000 929.200000 21.075000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.304 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.33 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.486 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.540000 0.000000 0.840000 0.800000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 67.220000 0.800000 67.520000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 134.585000 0.800000 134.885000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 201.955000 0.800000 202.255000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 269.320000 0.800000 269.620000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 336.690000 0.800000 336.990000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 404.060000 0.800000 404.360000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 471.425000 0.800000 471.725000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 538.795000 0.800000 539.095000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 606.160000 0.800000 606.460000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 673.530000 0.800000 673.830000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 740.900000 0.800000 741.200000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 808.265000 0.800000 808.565000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 875.635000 0.800000 875.935000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 129.459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 644.78 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.6 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 15.340000 920.230000 15.480000 920.720000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 129.435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 644.658 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.6 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 107.145000 920.230000 107.285000 920.720000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 129.459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 644.78 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.6 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 214.360000 920.230000 214.500000 920.720000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 129.435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 644.658 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.6 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 321.570000 920.230000 321.710000 920.720000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 129.435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 644.658 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.6 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 428.785000 920.230000 428.925000 920.720000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 129.459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 644.78 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.6 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 536.000000 920.230000 536.140000 920.720000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 129.459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 644.78 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.6 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 643.215000 920.230000 643.355000 920.720000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 129.459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 644.78 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.6 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 750.430000 920.230000 750.570000 920.720000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1382.76 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 129.425 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 644.511 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.6 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 173.669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 943.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 857.640000 920.230000 857.780000 920.720000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.37 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.68 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.531 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 911.190000 929.200000 911.490000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 857.775000 929.200000 858.075000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 795.000000 929.200000 795.300000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 732.225000 929.200000 732.525000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 669.450000 929.200000 669.750000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 606.675000 929.200000 606.975000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.37 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.68 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.531 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 543.900000 929.200000 544.200000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 481.125000 929.200000 481.425000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.37 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.68 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.531 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 418.350000 929.200000 418.650000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 119.066 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 635.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.7271 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 213.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 9.828 LAYER met4  ;
    ANTENNAMAXAREACAR 17.5338 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 84.64 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.332936 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 355.575000 929.200000 355.875000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 292.800000 929.200000 293.100000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.37 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.68 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.531 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 230.025000 929.200000 230.325000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.37 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.68 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.531 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 167.250000 929.200000 167.550000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.24 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 104.475000 929.200000 104.775000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.37 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.68 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.531 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.1148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.056 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 42.4509 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 69.3052 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 928.400000 41.700000 929.200000 42.000000 ;
    END
  END io_oeb[0]
  PIN irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.353 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1381.59 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.519 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 16.320000 0.800000 16.620000 ;
    END
  END irq[2]
  PIN irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 378.62 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1980.88 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.970623 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 173.519 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 44.6517 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 213.122 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 1.32243 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 87.1026 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 282.427 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 12.050000 0.800000 12.350000 ;
    END
  END irq[1]
  PIN irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met3  ;
    ANTENNAMAXAREACAR 254.221 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1380.18 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.429 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 941.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.224 LAYER met4  ;
    ANTENNAGATEAREA 0.6822 LAYER met4  ;
    ANTENNAMAXAREACAR 27.6294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.447 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.938141 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met5  ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 214.752 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 8.390000 0.800000 8.690000 ;
    END
  END irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 925.140000 2.100000 927.140000 918.620000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.060000 2.100000 4.060000 918.620000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 913.260000 511.650000 915.000000 906.430000 ;
      LAYER met4 ;
        RECT 437.940000 511.650000 439.680000 906.430000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 921.140000 6.100000 923.140000 914.620000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.060000 6.100000 8.060000 914.620000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 441.340000 515.050000 443.080000 903.030000 ;
      LAYER met4 ;
        RECT 909.860000 515.050000 911.600000 903.030000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 929.200000 920.720000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 929.200000 920.720000 ;
    LAYER met2 ;
      RECT 915.840000 920.090000 929.200000 920.720000 ;
      RECT 893.660000 920.090000 915.420000 920.720000 ;
      RECT 857.920000 920.090000 893.240000 920.720000 ;
      RECT 822.185000 920.090000 857.500000 920.720000 ;
      RECT 786.445000 920.090000 821.765000 920.720000 ;
      RECT 750.710000 920.090000 786.025000 920.720000 ;
      RECT 714.970000 920.090000 750.290000 920.720000 ;
      RECT 679.230000 920.090000 714.550000 920.720000 ;
      RECT 643.495000 920.090000 678.810000 920.720000 ;
      RECT 607.755000 920.090000 643.075000 920.720000 ;
      RECT 572.020000 920.090000 607.335000 920.720000 ;
      RECT 536.280000 920.090000 571.600000 920.720000 ;
      RECT 500.540000 920.090000 535.860000 920.720000 ;
      RECT 464.805000 920.090000 500.120000 920.720000 ;
      RECT 429.065000 920.090000 464.385000 920.720000 ;
      RECT 393.330000 920.090000 428.645000 920.720000 ;
      RECT 357.590000 920.090000 392.910000 920.720000 ;
      RECT 321.850000 920.090000 357.170000 920.720000 ;
      RECT 286.115000 920.090000 321.430000 920.720000 ;
      RECT 250.375000 920.090000 285.695000 920.720000 ;
      RECT 214.640000 920.090000 249.955000 920.720000 ;
      RECT 178.900000 920.090000 214.220000 920.720000 ;
      RECT 143.160000 920.090000 178.480000 920.720000 ;
      RECT 107.425000 920.090000 142.740000 920.720000 ;
      RECT 71.685000 920.090000 107.005000 920.720000 ;
      RECT 35.950000 920.090000 71.265000 920.720000 ;
      RECT 15.620000 920.090000 35.530000 920.720000 ;
      RECT 0.000000 920.090000 15.200000 920.720000 ;
      RECT 0.000000 4.460000 929.200000 920.090000 ;
      RECT 0.630000 4.040000 929.200000 4.460000 ;
      RECT 0.000000 0.630000 929.200000 4.040000 ;
      RECT 927.410000 0.000000 928.890000 0.630000 ;
      RECT 925.510000 0.000000 926.990000 0.630000 ;
      RECT 923.610000 0.000000 925.090000 0.630000 ;
      RECT 921.710000 0.000000 923.190000 0.630000 ;
      RECT 919.810000 0.000000 921.290000 0.630000 ;
      RECT 917.910000 0.000000 919.390000 0.630000 ;
      RECT 916.010000 0.000000 917.490000 0.630000 ;
      RECT 914.110000 0.000000 915.590000 0.630000 ;
      RECT 912.210000 0.000000 913.690000 0.630000 ;
      RECT 910.310000 0.000000 911.790000 0.630000 ;
      RECT 908.410000 0.000000 909.890000 0.630000 ;
      RECT 906.510000 0.000000 907.990000 0.630000 ;
      RECT 904.610000 0.000000 906.090000 0.630000 ;
      RECT 902.710000 0.000000 904.190000 0.630000 ;
      RECT 900.810000 0.000000 902.290000 0.630000 ;
      RECT 898.910000 0.000000 900.390000 0.630000 ;
      RECT 897.010000 0.000000 898.490000 0.630000 ;
      RECT 895.110000 0.000000 896.590000 0.630000 ;
      RECT 893.210000 0.000000 894.690000 0.630000 ;
      RECT 891.310000 0.000000 892.790000 0.630000 ;
      RECT 889.410000 0.000000 890.890000 0.630000 ;
      RECT 887.510000 0.000000 888.990000 0.630000 ;
      RECT 885.610000 0.000000 887.090000 0.630000 ;
      RECT 883.710000 0.000000 885.190000 0.630000 ;
      RECT 881.810000 0.000000 883.290000 0.630000 ;
      RECT 879.910000 0.000000 881.390000 0.630000 ;
      RECT 878.010000 0.000000 879.490000 0.630000 ;
      RECT 876.110000 0.000000 877.590000 0.630000 ;
      RECT 874.210000 0.000000 875.690000 0.630000 ;
      RECT 872.310000 0.000000 873.790000 0.630000 ;
      RECT 870.410000 0.000000 871.890000 0.630000 ;
      RECT 868.510000 0.000000 869.990000 0.630000 ;
      RECT 866.610000 0.000000 868.090000 0.630000 ;
      RECT 864.710000 0.000000 866.190000 0.630000 ;
      RECT 862.810000 0.000000 864.290000 0.630000 ;
      RECT 860.910000 0.000000 862.390000 0.630000 ;
      RECT 859.010000 0.000000 860.490000 0.630000 ;
      RECT 857.110000 0.000000 858.590000 0.630000 ;
      RECT 855.210000 0.000000 856.690000 0.630000 ;
      RECT 853.310000 0.000000 854.790000 0.630000 ;
      RECT 851.410000 0.000000 852.890000 0.630000 ;
      RECT 849.510000 0.000000 850.990000 0.630000 ;
      RECT 847.610000 0.000000 849.090000 0.630000 ;
      RECT 845.710000 0.000000 847.190000 0.630000 ;
      RECT 843.810000 0.000000 845.290000 0.630000 ;
      RECT 841.910000 0.000000 843.390000 0.630000 ;
      RECT 840.010000 0.000000 841.490000 0.630000 ;
      RECT 838.110000 0.000000 839.590000 0.630000 ;
      RECT 836.210000 0.000000 837.690000 0.630000 ;
      RECT 834.310000 0.000000 835.790000 0.630000 ;
      RECT 832.410000 0.000000 833.890000 0.630000 ;
      RECT 830.510000 0.000000 831.990000 0.630000 ;
      RECT 828.610000 0.000000 830.090000 0.630000 ;
      RECT 826.710000 0.000000 828.190000 0.630000 ;
      RECT 824.810000 0.000000 826.290000 0.630000 ;
      RECT 822.910000 0.000000 824.390000 0.630000 ;
      RECT 821.010000 0.000000 822.490000 0.630000 ;
      RECT 819.110000 0.000000 820.590000 0.630000 ;
      RECT 817.210000 0.000000 818.690000 0.630000 ;
      RECT 815.310000 0.000000 816.790000 0.630000 ;
      RECT 813.410000 0.000000 814.890000 0.630000 ;
      RECT 811.510000 0.000000 812.990000 0.630000 ;
      RECT 809.610000 0.000000 811.090000 0.630000 ;
      RECT 807.710000 0.000000 809.190000 0.630000 ;
      RECT 805.810000 0.000000 807.290000 0.630000 ;
      RECT 803.910000 0.000000 805.390000 0.630000 ;
      RECT 802.010000 0.000000 803.490000 0.630000 ;
      RECT 800.110000 0.000000 801.590000 0.630000 ;
      RECT 798.210000 0.000000 799.690000 0.630000 ;
      RECT 796.310000 0.000000 797.790000 0.630000 ;
      RECT 794.410000 0.000000 795.890000 0.630000 ;
      RECT 792.510000 0.000000 793.990000 0.630000 ;
      RECT 790.610000 0.000000 792.090000 0.630000 ;
      RECT 788.710000 0.000000 790.190000 0.630000 ;
      RECT 786.810000 0.000000 788.290000 0.630000 ;
      RECT 784.910000 0.000000 786.390000 0.630000 ;
      RECT 783.010000 0.000000 784.490000 0.630000 ;
      RECT 781.110000 0.000000 782.590000 0.630000 ;
      RECT 779.210000 0.000000 780.690000 0.630000 ;
      RECT 777.310000 0.000000 778.790000 0.630000 ;
      RECT 775.410000 0.000000 776.890000 0.630000 ;
      RECT 773.510000 0.000000 774.990000 0.630000 ;
      RECT 771.610000 0.000000 773.090000 0.630000 ;
      RECT 769.710000 0.000000 771.190000 0.630000 ;
      RECT 767.810000 0.000000 769.290000 0.630000 ;
      RECT 765.910000 0.000000 767.390000 0.630000 ;
      RECT 764.010000 0.000000 765.490000 0.630000 ;
      RECT 762.110000 0.000000 763.590000 0.630000 ;
      RECT 760.210000 0.000000 761.690000 0.630000 ;
      RECT 758.310000 0.000000 759.790000 0.630000 ;
      RECT 756.410000 0.000000 757.890000 0.630000 ;
      RECT 754.510000 0.000000 755.990000 0.630000 ;
      RECT 752.610000 0.000000 754.090000 0.630000 ;
      RECT 750.710000 0.000000 752.190000 0.630000 ;
      RECT 748.810000 0.000000 750.290000 0.630000 ;
      RECT 746.910000 0.000000 748.390000 0.630000 ;
      RECT 745.010000 0.000000 746.490000 0.630000 ;
      RECT 743.110000 0.000000 744.590000 0.630000 ;
      RECT 741.210000 0.000000 742.690000 0.630000 ;
      RECT 739.310000 0.000000 740.790000 0.630000 ;
      RECT 737.410000 0.000000 738.890000 0.630000 ;
      RECT 735.510000 0.000000 736.990000 0.630000 ;
      RECT 733.610000 0.000000 735.090000 0.630000 ;
      RECT 731.710000 0.000000 733.190000 0.630000 ;
      RECT 729.810000 0.000000 731.290000 0.630000 ;
      RECT 727.910000 0.000000 729.390000 0.630000 ;
      RECT 726.010000 0.000000 727.490000 0.630000 ;
      RECT 724.110000 0.000000 725.590000 0.630000 ;
      RECT 722.210000 0.000000 723.690000 0.630000 ;
      RECT 720.310000 0.000000 721.790000 0.630000 ;
      RECT 718.410000 0.000000 719.890000 0.630000 ;
      RECT 716.510000 0.000000 717.990000 0.630000 ;
      RECT 714.610000 0.000000 716.090000 0.630000 ;
      RECT 712.710000 0.000000 714.190000 0.630000 ;
      RECT 710.810000 0.000000 712.290000 0.630000 ;
      RECT 708.910000 0.000000 710.390000 0.630000 ;
      RECT 707.010000 0.000000 708.490000 0.630000 ;
      RECT 705.110000 0.000000 706.590000 0.630000 ;
      RECT 703.210000 0.000000 704.690000 0.630000 ;
      RECT 701.310000 0.000000 702.790000 0.630000 ;
      RECT 699.410000 0.000000 700.890000 0.630000 ;
      RECT 697.510000 0.000000 698.990000 0.630000 ;
      RECT 695.610000 0.000000 697.090000 0.630000 ;
      RECT 693.710000 0.000000 695.190000 0.630000 ;
      RECT 691.810000 0.000000 693.290000 0.630000 ;
      RECT 689.910000 0.000000 691.390000 0.630000 ;
      RECT 688.010000 0.000000 689.490000 0.630000 ;
      RECT 686.110000 0.000000 687.590000 0.630000 ;
      RECT 684.210000 0.000000 685.690000 0.630000 ;
      RECT 682.310000 0.000000 683.790000 0.630000 ;
      RECT 680.410000 0.000000 681.890000 0.630000 ;
      RECT 678.510000 0.000000 679.990000 0.630000 ;
      RECT 676.610000 0.000000 678.090000 0.630000 ;
      RECT 674.710000 0.000000 676.190000 0.630000 ;
      RECT 672.810000 0.000000 674.290000 0.630000 ;
      RECT 670.910000 0.000000 672.390000 0.630000 ;
      RECT 669.010000 0.000000 670.490000 0.630000 ;
      RECT 667.110000 0.000000 668.590000 0.630000 ;
      RECT 665.210000 0.000000 666.690000 0.630000 ;
      RECT 663.310000 0.000000 664.790000 0.630000 ;
      RECT 661.410000 0.000000 662.890000 0.630000 ;
      RECT 659.510000 0.000000 660.990000 0.630000 ;
      RECT 657.610000 0.000000 659.090000 0.630000 ;
      RECT 655.710000 0.000000 657.190000 0.630000 ;
      RECT 653.810000 0.000000 655.290000 0.630000 ;
      RECT 651.910000 0.000000 653.390000 0.630000 ;
      RECT 650.010000 0.000000 651.490000 0.630000 ;
      RECT 648.110000 0.000000 649.590000 0.630000 ;
      RECT 646.210000 0.000000 647.690000 0.630000 ;
      RECT 644.310000 0.000000 645.790000 0.630000 ;
      RECT 642.410000 0.000000 643.890000 0.630000 ;
      RECT 640.510000 0.000000 641.990000 0.630000 ;
      RECT 638.610000 0.000000 640.090000 0.630000 ;
      RECT 636.710000 0.000000 638.190000 0.630000 ;
      RECT 634.810000 0.000000 636.290000 0.630000 ;
      RECT 632.910000 0.000000 634.390000 0.630000 ;
      RECT 631.010000 0.000000 632.490000 0.630000 ;
      RECT 629.110000 0.000000 630.590000 0.630000 ;
      RECT 627.210000 0.000000 628.690000 0.630000 ;
      RECT 625.310000 0.000000 626.790000 0.630000 ;
      RECT 623.410000 0.000000 624.890000 0.630000 ;
      RECT 621.510000 0.000000 622.990000 0.630000 ;
      RECT 619.610000 0.000000 621.090000 0.630000 ;
      RECT 617.710000 0.000000 619.190000 0.630000 ;
      RECT 615.810000 0.000000 617.290000 0.630000 ;
      RECT 613.910000 0.000000 615.390000 0.630000 ;
      RECT 612.010000 0.000000 613.490000 0.630000 ;
      RECT 610.110000 0.000000 611.590000 0.630000 ;
      RECT 608.210000 0.000000 609.690000 0.630000 ;
      RECT 606.310000 0.000000 607.790000 0.630000 ;
      RECT 604.410000 0.000000 605.890000 0.630000 ;
      RECT 602.510000 0.000000 603.990000 0.630000 ;
      RECT 600.610000 0.000000 602.090000 0.630000 ;
      RECT 598.710000 0.000000 600.190000 0.630000 ;
      RECT 596.810000 0.000000 598.290000 0.630000 ;
      RECT 594.910000 0.000000 596.390000 0.630000 ;
      RECT 593.010000 0.000000 594.490000 0.630000 ;
      RECT 591.110000 0.000000 592.590000 0.630000 ;
      RECT 589.210000 0.000000 590.690000 0.630000 ;
      RECT 587.310000 0.000000 588.790000 0.630000 ;
      RECT 585.410000 0.000000 586.890000 0.630000 ;
      RECT 583.510000 0.000000 584.990000 0.630000 ;
      RECT 581.610000 0.000000 583.090000 0.630000 ;
      RECT 579.710000 0.000000 581.190000 0.630000 ;
      RECT 577.810000 0.000000 579.290000 0.630000 ;
      RECT 575.910000 0.000000 577.390000 0.630000 ;
      RECT 574.010000 0.000000 575.490000 0.630000 ;
      RECT 572.110000 0.000000 573.590000 0.630000 ;
      RECT 570.210000 0.000000 571.690000 0.630000 ;
      RECT 568.310000 0.000000 569.790000 0.630000 ;
      RECT 566.410000 0.000000 567.890000 0.630000 ;
      RECT 564.510000 0.000000 565.990000 0.630000 ;
      RECT 562.610000 0.000000 564.090000 0.630000 ;
      RECT 560.710000 0.000000 562.190000 0.630000 ;
      RECT 558.810000 0.000000 560.290000 0.630000 ;
      RECT 556.910000 0.000000 558.390000 0.630000 ;
      RECT 555.010000 0.000000 556.490000 0.630000 ;
      RECT 553.110000 0.000000 554.590000 0.630000 ;
      RECT 551.210000 0.000000 552.690000 0.630000 ;
      RECT 549.310000 0.000000 550.790000 0.630000 ;
      RECT 547.410000 0.000000 548.890000 0.630000 ;
      RECT 545.510000 0.000000 546.990000 0.630000 ;
      RECT 543.610000 0.000000 545.090000 0.630000 ;
      RECT 541.710000 0.000000 543.190000 0.630000 ;
      RECT 539.810000 0.000000 541.290000 0.630000 ;
      RECT 537.910000 0.000000 539.390000 0.630000 ;
      RECT 536.010000 0.000000 537.490000 0.630000 ;
      RECT 534.110000 0.000000 535.590000 0.630000 ;
      RECT 532.210000 0.000000 533.690000 0.630000 ;
      RECT 530.310000 0.000000 531.790000 0.630000 ;
      RECT 528.410000 0.000000 529.890000 0.630000 ;
      RECT 526.510000 0.000000 527.990000 0.630000 ;
      RECT 524.610000 0.000000 526.090000 0.630000 ;
      RECT 522.710000 0.000000 524.190000 0.630000 ;
      RECT 520.810000 0.000000 522.290000 0.630000 ;
      RECT 518.910000 0.000000 520.390000 0.630000 ;
      RECT 517.010000 0.000000 518.490000 0.630000 ;
      RECT 515.110000 0.000000 516.590000 0.630000 ;
      RECT 513.210000 0.000000 514.690000 0.630000 ;
      RECT 511.310000 0.000000 512.790000 0.630000 ;
      RECT 509.410000 0.000000 510.890000 0.630000 ;
      RECT 507.510000 0.000000 508.990000 0.630000 ;
      RECT 505.610000 0.000000 507.090000 0.630000 ;
      RECT 503.710000 0.000000 505.190000 0.630000 ;
      RECT 501.810000 0.000000 503.290000 0.630000 ;
      RECT 499.910000 0.000000 501.390000 0.630000 ;
      RECT 498.010000 0.000000 499.490000 0.630000 ;
      RECT 496.110000 0.000000 497.590000 0.630000 ;
      RECT 494.210000 0.000000 495.690000 0.630000 ;
      RECT 492.310000 0.000000 493.790000 0.630000 ;
      RECT 490.410000 0.000000 491.890000 0.630000 ;
      RECT 488.510000 0.000000 489.990000 0.630000 ;
      RECT 486.610000 0.000000 488.090000 0.630000 ;
      RECT 484.710000 0.000000 486.190000 0.630000 ;
      RECT 482.810000 0.000000 484.290000 0.630000 ;
      RECT 480.910000 0.000000 482.390000 0.630000 ;
      RECT 479.010000 0.000000 480.490000 0.630000 ;
      RECT 477.110000 0.000000 478.590000 0.630000 ;
      RECT 475.210000 0.000000 476.690000 0.630000 ;
      RECT 473.310000 0.000000 474.790000 0.630000 ;
      RECT 471.410000 0.000000 472.890000 0.630000 ;
      RECT 469.510000 0.000000 470.990000 0.630000 ;
      RECT 467.610000 0.000000 469.090000 0.630000 ;
      RECT 465.710000 0.000000 467.190000 0.630000 ;
      RECT 463.810000 0.000000 465.290000 0.630000 ;
      RECT 461.910000 0.000000 463.390000 0.630000 ;
      RECT 460.010000 0.000000 461.490000 0.630000 ;
      RECT 458.110000 0.000000 459.590000 0.630000 ;
      RECT 456.210000 0.000000 457.690000 0.630000 ;
      RECT 454.310000 0.000000 455.790000 0.630000 ;
      RECT 452.410000 0.000000 453.890000 0.630000 ;
      RECT 450.510000 0.000000 451.990000 0.630000 ;
      RECT 448.610000 0.000000 450.090000 0.630000 ;
      RECT 446.710000 0.000000 448.190000 0.630000 ;
      RECT 444.810000 0.000000 446.290000 0.630000 ;
      RECT 442.910000 0.000000 444.390000 0.630000 ;
      RECT 441.010000 0.000000 442.490000 0.630000 ;
      RECT 439.110000 0.000000 440.590000 0.630000 ;
      RECT 437.210000 0.000000 438.690000 0.630000 ;
      RECT 435.310000 0.000000 436.790000 0.630000 ;
      RECT 433.410000 0.000000 434.890000 0.630000 ;
      RECT 431.510000 0.000000 432.990000 0.630000 ;
      RECT 429.610000 0.000000 431.090000 0.630000 ;
      RECT 427.710000 0.000000 429.190000 0.630000 ;
      RECT 425.810000 0.000000 427.290000 0.630000 ;
      RECT 423.910000 0.000000 425.390000 0.630000 ;
      RECT 422.010000 0.000000 423.490000 0.630000 ;
      RECT 420.110000 0.000000 421.590000 0.630000 ;
      RECT 418.210000 0.000000 419.690000 0.630000 ;
      RECT 416.310000 0.000000 417.790000 0.630000 ;
      RECT 414.410000 0.000000 415.890000 0.630000 ;
      RECT 412.510000 0.000000 413.990000 0.630000 ;
      RECT 410.610000 0.000000 412.090000 0.630000 ;
      RECT 408.710000 0.000000 410.190000 0.630000 ;
      RECT 406.810000 0.000000 408.290000 0.630000 ;
      RECT 404.910000 0.000000 406.390000 0.630000 ;
      RECT 403.010000 0.000000 404.490000 0.630000 ;
      RECT 401.110000 0.000000 402.590000 0.630000 ;
      RECT 399.210000 0.000000 400.690000 0.630000 ;
      RECT 397.310000 0.000000 398.790000 0.630000 ;
      RECT 395.410000 0.000000 396.890000 0.630000 ;
      RECT 393.510000 0.000000 394.990000 0.630000 ;
      RECT 391.610000 0.000000 393.090000 0.630000 ;
      RECT 389.710000 0.000000 391.190000 0.630000 ;
      RECT 387.810000 0.000000 389.290000 0.630000 ;
      RECT 385.910000 0.000000 387.390000 0.630000 ;
      RECT 384.010000 0.000000 385.490000 0.630000 ;
      RECT 382.110000 0.000000 383.590000 0.630000 ;
      RECT 380.210000 0.000000 381.690000 0.630000 ;
      RECT 378.310000 0.000000 379.790000 0.630000 ;
      RECT 376.410000 0.000000 377.890000 0.630000 ;
      RECT 374.510000 0.000000 375.990000 0.630000 ;
      RECT 372.610000 0.000000 374.090000 0.630000 ;
      RECT 370.710000 0.000000 372.190000 0.630000 ;
      RECT 368.810000 0.000000 370.290000 0.630000 ;
      RECT 366.910000 0.000000 368.390000 0.630000 ;
      RECT 365.010000 0.000000 366.490000 0.630000 ;
      RECT 363.110000 0.000000 364.590000 0.630000 ;
      RECT 361.210000 0.000000 362.690000 0.630000 ;
      RECT 359.310000 0.000000 360.790000 0.630000 ;
      RECT 357.410000 0.000000 358.890000 0.630000 ;
      RECT 355.510000 0.000000 356.990000 0.630000 ;
      RECT 353.610000 0.000000 355.090000 0.630000 ;
      RECT 351.710000 0.000000 353.190000 0.630000 ;
      RECT 349.810000 0.000000 351.290000 0.630000 ;
      RECT 347.910000 0.000000 349.390000 0.630000 ;
      RECT 346.010000 0.000000 347.490000 0.630000 ;
      RECT 344.110000 0.000000 345.590000 0.630000 ;
      RECT 342.210000 0.000000 343.690000 0.630000 ;
      RECT 340.310000 0.000000 341.790000 0.630000 ;
      RECT 338.410000 0.000000 339.890000 0.630000 ;
      RECT 336.510000 0.000000 337.990000 0.630000 ;
      RECT 334.610000 0.000000 336.090000 0.630000 ;
      RECT 332.710000 0.000000 334.190000 0.630000 ;
      RECT 330.810000 0.000000 332.290000 0.630000 ;
      RECT 328.910000 0.000000 330.390000 0.630000 ;
      RECT 327.010000 0.000000 328.490000 0.630000 ;
      RECT 325.110000 0.000000 326.590000 0.630000 ;
      RECT 323.210000 0.000000 324.690000 0.630000 ;
      RECT 321.310000 0.000000 322.790000 0.630000 ;
      RECT 319.410000 0.000000 320.890000 0.630000 ;
      RECT 317.510000 0.000000 318.990000 0.630000 ;
      RECT 315.610000 0.000000 317.090000 0.630000 ;
      RECT 313.710000 0.000000 315.190000 0.630000 ;
      RECT 311.810000 0.000000 313.290000 0.630000 ;
      RECT 309.910000 0.000000 311.390000 0.630000 ;
      RECT 308.010000 0.000000 309.490000 0.630000 ;
      RECT 306.110000 0.000000 307.590000 0.630000 ;
      RECT 304.210000 0.000000 305.690000 0.630000 ;
      RECT 302.310000 0.000000 303.790000 0.630000 ;
      RECT 300.410000 0.000000 301.890000 0.630000 ;
      RECT 298.510000 0.000000 299.990000 0.630000 ;
      RECT 296.610000 0.000000 298.090000 0.630000 ;
      RECT 294.710000 0.000000 296.190000 0.630000 ;
      RECT 292.810000 0.000000 294.290000 0.630000 ;
      RECT 290.910000 0.000000 292.390000 0.630000 ;
      RECT 289.010000 0.000000 290.490000 0.630000 ;
      RECT 287.110000 0.000000 288.590000 0.630000 ;
      RECT 285.210000 0.000000 286.690000 0.630000 ;
      RECT 283.310000 0.000000 284.790000 0.630000 ;
      RECT 281.410000 0.000000 282.890000 0.630000 ;
      RECT 279.510000 0.000000 280.990000 0.630000 ;
      RECT 277.610000 0.000000 279.090000 0.630000 ;
      RECT 275.710000 0.000000 277.190000 0.630000 ;
      RECT 273.810000 0.000000 275.290000 0.630000 ;
      RECT 271.910000 0.000000 273.390000 0.630000 ;
      RECT 270.010000 0.000000 271.490000 0.630000 ;
      RECT 268.110000 0.000000 269.590000 0.630000 ;
      RECT 266.210000 0.000000 267.690000 0.630000 ;
      RECT 264.310000 0.000000 265.790000 0.630000 ;
      RECT 262.410000 0.000000 263.890000 0.630000 ;
      RECT 260.510000 0.000000 261.990000 0.630000 ;
      RECT 258.610000 0.000000 260.090000 0.630000 ;
      RECT 256.710000 0.000000 258.190000 0.630000 ;
      RECT 254.810000 0.000000 256.290000 0.630000 ;
      RECT 252.910000 0.000000 254.390000 0.630000 ;
      RECT 251.010000 0.000000 252.490000 0.630000 ;
      RECT 249.110000 0.000000 250.590000 0.630000 ;
      RECT 247.210000 0.000000 248.690000 0.630000 ;
      RECT 245.310000 0.000000 246.790000 0.630000 ;
      RECT 243.410000 0.000000 244.890000 0.630000 ;
      RECT 241.510000 0.000000 242.990000 0.630000 ;
      RECT 239.610000 0.000000 241.090000 0.630000 ;
      RECT 237.710000 0.000000 239.190000 0.630000 ;
      RECT 235.810000 0.000000 237.290000 0.630000 ;
      RECT 233.910000 0.000000 235.390000 0.630000 ;
      RECT 232.010000 0.000000 233.490000 0.630000 ;
      RECT 230.110000 0.000000 231.590000 0.630000 ;
      RECT 228.210000 0.000000 229.690000 0.630000 ;
      RECT 226.310000 0.000000 227.790000 0.630000 ;
      RECT 224.410000 0.000000 225.890000 0.630000 ;
      RECT 222.510000 0.000000 223.990000 0.630000 ;
      RECT 220.610000 0.000000 222.090000 0.630000 ;
      RECT 218.710000 0.000000 220.190000 0.630000 ;
      RECT 216.810000 0.000000 218.290000 0.630000 ;
      RECT 214.910000 0.000000 216.390000 0.630000 ;
      RECT 213.010000 0.000000 214.490000 0.630000 ;
      RECT 211.110000 0.000000 212.590000 0.630000 ;
      RECT 209.210000 0.000000 210.690000 0.630000 ;
      RECT 207.310000 0.000000 208.790000 0.630000 ;
      RECT 205.410000 0.000000 206.890000 0.630000 ;
      RECT 203.510000 0.000000 204.990000 0.630000 ;
      RECT 201.610000 0.000000 203.090000 0.630000 ;
      RECT 199.710000 0.000000 201.190000 0.630000 ;
      RECT 197.810000 0.000000 199.290000 0.630000 ;
      RECT 195.910000 0.000000 197.390000 0.630000 ;
      RECT 194.010000 0.000000 195.490000 0.630000 ;
      RECT 192.110000 0.000000 193.590000 0.630000 ;
      RECT 190.210000 0.000000 191.690000 0.630000 ;
      RECT 188.310000 0.000000 189.790000 0.630000 ;
      RECT 186.410000 0.000000 187.890000 0.630000 ;
      RECT 184.510000 0.000000 185.990000 0.630000 ;
      RECT 182.610000 0.000000 184.090000 0.630000 ;
      RECT 180.710000 0.000000 182.190000 0.630000 ;
      RECT 178.810000 0.000000 180.290000 0.630000 ;
      RECT 176.910000 0.000000 178.390000 0.630000 ;
      RECT 175.010000 0.000000 176.490000 0.630000 ;
      RECT 173.110000 0.000000 174.590000 0.630000 ;
      RECT 171.210000 0.000000 172.690000 0.630000 ;
      RECT 169.310000 0.000000 170.790000 0.630000 ;
      RECT 167.410000 0.000000 168.890000 0.630000 ;
      RECT 165.510000 0.000000 166.990000 0.630000 ;
      RECT 163.610000 0.000000 165.090000 0.630000 ;
      RECT 161.710000 0.000000 163.190000 0.630000 ;
      RECT 159.810000 0.000000 161.290000 0.630000 ;
      RECT 157.910000 0.000000 159.390000 0.630000 ;
      RECT 156.010000 0.000000 157.490000 0.630000 ;
      RECT 154.110000 0.000000 155.590000 0.630000 ;
      RECT 152.210000 0.000000 153.690000 0.630000 ;
      RECT 150.310000 0.000000 151.790000 0.630000 ;
      RECT 148.410000 0.000000 149.890000 0.630000 ;
      RECT 146.510000 0.000000 147.990000 0.630000 ;
      RECT 144.610000 0.000000 146.090000 0.630000 ;
      RECT 142.710000 0.000000 144.190000 0.630000 ;
      RECT 140.810000 0.000000 142.290000 0.630000 ;
      RECT 138.910000 0.000000 140.390000 0.630000 ;
      RECT 137.010000 0.000000 138.490000 0.630000 ;
      RECT 135.110000 0.000000 136.590000 0.630000 ;
      RECT 133.210000 0.000000 134.690000 0.630000 ;
      RECT 131.310000 0.000000 132.790000 0.630000 ;
      RECT 129.410000 0.000000 130.890000 0.630000 ;
      RECT 127.510000 0.000000 128.990000 0.630000 ;
      RECT 125.610000 0.000000 127.090000 0.630000 ;
      RECT 123.710000 0.000000 125.190000 0.630000 ;
      RECT 121.810000 0.000000 123.290000 0.630000 ;
      RECT 119.910000 0.000000 121.390000 0.630000 ;
      RECT 118.010000 0.000000 119.490000 0.630000 ;
      RECT 116.110000 0.000000 117.590000 0.630000 ;
      RECT 114.210000 0.000000 115.690000 0.630000 ;
      RECT 112.310000 0.000000 113.790000 0.630000 ;
      RECT 110.410000 0.000000 111.890000 0.630000 ;
      RECT 108.510000 0.000000 109.990000 0.630000 ;
      RECT 106.610000 0.000000 108.090000 0.630000 ;
      RECT 104.710000 0.000000 106.190000 0.630000 ;
      RECT 102.810000 0.000000 104.290000 0.630000 ;
      RECT 100.910000 0.000000 102.390000 0.630000 ;
      RECT 99.010000 0.000000 100.490000 0.630000 ;
      RECT 97.110000 0.000000 98.590000 0.630000 ;
      RECT 95.210000 0.000000 96.690000 0.630000 ;
      RECT 93.310000 0.000000 94.790000 0.630000 ;
      RECT 91.410000 0.000000 92.890000 0.630000 ;
      RECT 89.510000 0.000000 90.990000 0.630000 ;
      RECT 87.610000 0.000000 89.090000 0.630000 ;
      RECT 85.710000 0.000000 87.190000 0.630000 ;
      RECT 83.810000 0.000000 85.290000 0.630000 ;
      RECT 81.910000 0.000000 83.390000 0.630000 ;
      RECT 80.010000 0.000000 81.490000 0.630000 ;
      RECT 78.110000 0.000000 79.590000 0.630000 ;
      RECT 76.210000 0.000000 77.690000 0.630000 ;
      RECT 74.310000 0.000000 75.790000 0.630000 ;
      RECT 72.410000 0.000000 73.890000 0.630000 ;
      RECT 70.510000 0.000000 71.990000 0.630000 ;
      RECT 68.610000 0.000000 70.090000 0.630000 ;
      RECT 66.710000 0.000000 68.190000 0.630000 ;
      RECT 64.810000 0.000000 66.290000 0.630000 ;
      RECT 62.910000 0.000000 64.390000 0.630000 ;
      RECT 61.010000 0.000000 62.490000 0.630000 ;
      RECT 59.110000 0.000000 60.590000 0.630000 ;
      RECT 57.210000 0.000000 58.690000 0.630000 ;
      RECT 55.310000 0.000000 56.790000 0.630000 ;
      RECT 53.410000 0.000000 54.890000 0.630000 ;
      RECT 51.510000 0.000000 52.990000 0.630000 ;
      RECT 49.610000 0.000000 51.090000 0.630000 ;
      RECT 47.710000 0.000000 49.190000 0.630000 ;
      RECT 45.810000 0.000000 47.290000 0.630000 ;
      RECT 43.910000 0.000000 45.390000 0.630000 ;
      RECT 42.010000 0.000000 43.490000 0.630000 ;
      RECT 40.110000 0.000000 41.590000 0.630000 ;
      RECT 38.210000 0.000000 39.690000 0.630000 ;
      RECT 36.310000 0.000000 37.790000 0.630000 ;
      RECT 34.410000 0.000000 35.890000 0.630000 ;
      RECT 32.510000 0.000000 33.990000 0.630000 ;
      RECT 30.610000 0.000000 32.090000 0.630000 ;
      RECT 28.710000 0.000000 30.190000 0.630000 ;
      RECT 26.810000 0.000000 28.290000 0.630000 ;
      RECT 24.910000 0.000000 26.390000 0.630000 ;
      RECT 23.010000 0.000000 24.490000 0.630000 ;
      RECT 21.110000 0.000000 22.590000 0.630000 ;
      RECT 19.210000 0.000000 20.690000 0.630000 ;
      RECT 17.310000 0.000000 18.790000 0.630000 ;
      RECT 15.410000 0.000000 16.890000 0.630000 ;
      RECT 13.510000 0.000000 14.990000 0.630000 ;
      RECT 11.610000 0.000000 13.090000 0.630000 ;
      RECT 9.710000 0.000000 11.190000 0.630000 ;
      RECT 7.810000 0.000000 9.290000 0.630000 ;
      RECT 5.910000 0.000000 7.390000 0.630000 ;
      RECT 4.010000 0.000000 5.490000 0.630000 ;
      RECT 2.110000 0.000000 3.590000 0.630000 ;
      RECT 0.000000 0.000000 1.690000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 913.620000 929.200000 920.720000 ;
      RECT 1.100000 912.720000 929.200000 913.620000 ;
      RECT 0.000000 911.790000 929.200000 912.720000 ;
      RECT 0.000000 910.890000 928.100000 911.790000 ;
      RECT 0.000000 900.225000 929.200000 910.890000 ;
      RECT 0.000000 899.325000 928.100000 900.225000 ;
      RECT 0.000000 898.690000 929.200000 899.325000 ;
      RECT 1.100000 897.790000 929.200000 898.690000 ;
      RECT 0.000000 879.300000 929.200000 897.790000 ;
      RECT 0.000000 878.400000 928.100000 879.300000 ;
      RECT 0.000000 876.235000 929.200000 878.400000 ;
      RECT 1.100000 875.335000 929.200000 876.235000 ;
      RECT 0.000000 858.375000 929.200000 875.335000 ;
      RECT 0.000000 857.475000 928.100000 858.375000 ;
      RECT 0.000000 853.780000 929.200000 857.475000 ;
      RECT 1.100000 852.880000 929.200000 853.780000 ;
      RECT 0.000000 837.450000 929.200000 852.880000 ;
      RECT 0.000000 836.550000 928.100000 837.450000 ;
      RECT 0.000000 831.320000 929.200000 836.550000 ;
      RECT 1.100000 830.420000 929.200000 831.320000 ;
      RECT 0.000000 816.525000 929.200000 830.420000 ;
      RECT 0.000000 815.625000 928.100000 816.525000 ;
      RECT 0.000000 808.865000 929.200000 815.625000 ;
      RECT 1.100000 807.965000 929.200000 808.865000 ;
      RECT 0.000000 795.600000 929.200000 807.965000 ;
      RECT 0.000000 794.700000 928.100000 795.600000 ;
      RECT 0.000000 786.410000 929.200000 794.700000 ;
      RECT 1.100000 785.510000 929.200000 786.410000 ;
      RECT 0.000000 774.675000 929.200000 785.510000 ;
      RECT 0.000000 773.775000 928.100000 774.675000 ;
      RECT 0.000000 763.955000 929.200000 773.775000 ;
      RECT 1.100000 763.055000 929.200000 763.955000 ;
      RECT 0.000000 753.750000 929.200000 763.055000 ;
      RECT 0.000000 752.850000 928.100000 753.750000 ;
      RECT 0.000000 741.500000 929.200000 752.850000 ;
      RECT 1.100000 740.600000 929.200000 741.500000 ;
      RECT 0.000000 732.825000 929.200000 740.600000 ;
      RECT 0.000000 731.925000 928.100000 732.825000 ;
      RECT 0.000000 719.040000 929.200000 731.925000 ;
      RECT 1.100000 718.140000 929.200000 719.040000 ;
      RECT 0.000000 711.900000 929.200000 718.140000 ;
      RECT 0.000000 711.000000 928.100000 711.900000 ;
      RECT 0.000000 696.585000 929.200000 711.000000 ;
      RECT 1.100000 695.685000 929.200000 696.585000 ;
      RECT 0.000000 690.975000 929.200000 695.685000 ;
      RECT 0.000000 690.075000 928.100000 690.975000 ;
      RECT 0.000000 674.130000 929.200000 690.075000 ;
      RECT 1.100000 673.230000 929.200000 674.130000 ;
      RECT 0.000000 670.050000 929.200000 673.230000 ;
      RECT 0.000000 669.150000 928.100000 670.050000 ;
      RECT 0.000000 651.675000 929.200000 669.150000 ;
      RECT 1.100000 650.775000 929.200000 651.675000 ;
      RECT 0.000000 649.125000 929.200000 650.775000 ;
      RECT 0.000000 648.225000 928.100000 649.125000 ;
      RECT 0.000000 629.220000 929.200000 648.225000 ;
      RECT 1.100000 628.320000 929.200000 629.220000 ;
      RECT 0.000000 628.200000 929.200000 628.320000 ;
      RECT 0.000000 627.300000 928.100000 628.200000 ;
      RECT 0.000000 607.275000 929.200000 627.300000 ;
      RECT 0.000000 606.760000 928.100000 607.275000 ;
      RECT 1.100000 606.375000 928.100000 606.760000 ;
      RECT 1.100000 605.860000 929.200000 606.375000 ;
      RECT 0.000000 586.350000 929.200000 605.860000 ;
      RECT 0.000000 585.450000 928.100000 586.350000 ;
      RECT 0.000000 584.305000 929.200000 585.450000 ;
      RECT 1.100000 583.405000 929.200000 584.305000 ;
      RECT 0.000000 565.425000 929.200000 583.405000 ;
      RECT 0.000000 564.525000 928.100000 565.425000 ;
      RECT 0.000000 561.850000 929.200000 564.525000 ;
      RECT 1.100000 560.950000 929.200000 561.850000 ;
      RECT 0.000000 544.500000 929.200000 560.950000 ;
      RECT 0.000000 543.600000 928.100000 544.500000 ;
      RECT 0.000000 539.395000 929.200000 543.600000 ;
      RECT 1.100000 538.495000 929.200000 539.395000 ;
      RECT 0.000000 523.575000 929.200000 538.495000 ;
      RECT 0.000000 522.675000 928.100000 523.575000 ;
      RECT 0.000000 516.940000 929.200000 522.675000 ;
      RECT 1.100000 516.040000 929.200000 516.940000 ;
      RECT 0.000000 502.650000 929.200000 516.040000 ;
      RECT 0.000000 501.750000 928.100000 502.650000 ;
      RECT 0.000000 494.480000 929.200000 501.750000 ;
      RECT 1.100000 493.580000 929.200000 494.480000 ;
      RECT 0.000000 481.725000 929.200000 493.580000 ;
      RECT 0.000000 480.825000 928.100000 481.725000 ;
      RECT 0.000000 472.025000 929.200000 480.825000 ;
      RECT 1.100000 471.125000 929.200000 472.025000 ;
      RECT 0.000000 460.800000 929.200000 471.125000 ;
      RECT 0.000000 459.900000 928.100000 460.800000 ;
      RECT 0.000000 449.570000 929.200000 459.900000 ;
      RECT 1.100000 448.670000 929.200000 449.570000 ;
      RECT 0.000000 439.875000 929.200000 448.670000 ;
      RECT 0.000000 438.975000 928.100000 439.875000 ;
      RECT 0.000000 427.115000 929.200000 438.975000 ;
      RECT 1.100000 426.215000 929.200000 427.115000 ;
      RECT 0.000000 418.950000 929.200000 426.215000 ;
      RECT 0.000000 418.050000 928.100000 418.950000 ;
      RECT 0.000000 404.660000 929.200000 418.050000 ;
      RECT 1.100000 403.760000 929.200000 404.660000 ;
      RECT 0.000000 398.025000 929.200000 403.760000 ;
      RECT 0.000000 397.125000 928.100000 398.025000 ;
      RECT 0.000000 382.200000 929.200000 397.125000 ;
      RECT 1.100000 381.300000 929.200000 382.200000 ;
      RECT 0.000000 377.100000 929.200000 381.300000 ;
      RECT 0.000000 376.200000 928.100000 377.100000 ;
      RECT 0.000000 359.745000 929.200000 376.200000 ;
      RECT 1.100000 358.845000 929.200000 359.745000 ;
      RECT 0.000000 356.175000 929.200000 358.845000 ;
      RECT 0.000000 355.275000 928.100000 356.175000 ;
      RECT 0.000000 337.290000 929.200000 355.275000 ;
      RECT 1.100000 336.390000 929.200000 337.290000 ;
      RECT 0.000000 335.250000 929.200000 336.390000 ;
      RECT 0.000000 334.350000 928.100000 335.250000 ;
      RECT 0.000000 314.835000 929.200000 334.350000 ;
      RECT 1.100000 314.325000 929.200000 314.835000 ;
      RECT 1.100000 313.935000 928.100000 314.325000 ;
      RECT 0.000000 313.425000 928.100000 313.935000 ;
      RECT 0.000000 293.400000 929.200000 313.425000 ;
      RECT 0.000000 292.500000 928.100000 293.400000 ;
      RECT 0.000000 292.380000 929.200000 292.500000 ;
      RECT 1.100000 291.480000 929.200000 292.380000 ;
      RECT 0.000000 272.475000 929.200000 291.480000 ;
      RECT 0.000000 271.575000 928.100000 272.475000 ;
      RECT 0.000000 269.920000 929.200000 271.575000 ;
      RECT 1.100000 269.020000 929.200000 269.920000 ;
      RECT 0.000000 251.550000 929.200000 269.020000 ;
      RECT 0.000000 250.650000 928.100000 251.550000 ;
      RECT 0.000000 247.465000 929.200000 250.650000 ;
      RECT 1.100000 246.565000 929.200000 247.465000 ;
      RECT 0.000000 230.625000 929.200000 246.565000 ;
      RECT 0.000000 229.725000 928.100000 230.625000 ;
      RECT 0.000000 225.010000 929.200000 229.725000 ;
      RECT 1.100000 224.110000 929.200000 225.010000 ;
      RECT 0.000000 209.700000 929.200000 224.110000 ;
      RECT 0.000000 208.800000 928.100000 209.700000 ;
      RECT 0.000000 202.555000 929.200000 208.800000 ;
      RECT 1.100000 201.655000 929.200000 202.555000 ;
      RECT 0.000000 188.775000 929.200000 201.655000 ;
      RECT 0.000000 187.875000 928.100000 188.775000 ;
      RECT 0.000000 180.100000 929.200000 187.875000 ;
      RECT 1.100000 179.200000 929.200000 180.100000 ;
      RECT 0.000000 167.850000 929.200000 179.200000 ;
      RECT 0.000000 166.950000 928.100000 167.850000 ;
      RECT 0.000000 157.640000 929.200000 166.950000 ;
      RECT 1.100000 156.740000 929.200000 157.640000 ;
      RECT 0.000000 146.925000 929.200000 156.740000 ;
      RECT 0.000000 146.025000 928.100000 146.925000 ;
      RECT 0.000000 135.185000 929.200000 146.025000 ;
      RECT 1.100000 134.285000 929.200000 135.185000 ;
      RECT 0.000000 126.000000 929.200000 134.285000 ;
      RECT 0.000000 125.100000 928.100000 126.000000 ;
      RECT 0.000000 112.730000 929.200000 125.100000 ;
      RECT 1.100000 111.830000 929.200000 112.730000 ;
      RECT 0.000000 105.075000 929.200000 111.830000 ;
      RECT 0.000000 104.175000 928.100000 105.075000 ;
      RECT 0.000000 90.275000 929.200000 104.175000 ;
      RECT 1.100000 89.375000 929.200000 90.275000 ;
      RECT 0.000000 84.150000 929.200000 89.375000 ;
      RECT 0.000000 83.250000 928.100000 84.150000 ;
      RECT 0.000000 67.820000 929.200000 83.250000 ;
      RECT 1.100000 66.920000 929.200000 67.820000 ;
      RECT 0.000000 63.225000 929.200000 66.920000 ;
      RECT 0.000000 62.325000 928.100000 63.225000 ;
      RECT 0.000000 45.360000 929.200000 62.325000 ;
      RECT 1.100000 44.460000 929.200000 45.360000 ;
      RECT 0.000000 42.300000 929.200000 44.460000 ;
      RECT 0.000000 41.400000 928.100000 42.300000 ;
      RECT 0.000000 22.905000 929.200000 41.400000 ;
      RECT 1.100000 22.005000 929.200000 22.905000 ;
      RECT 0.000000 21.375000 929.200000 22.005000 ;
      RECT 0.000000 20.475000 928.100000 21.375000 ;
      RECT 0.000000 16.920000 929.200000 20.475000 ;
      RECT 1.100000 16.020000 929.200000 16.920000 ;
      RECT 0.000000 12.650000 929.200000 16.020000 ;
      RECT 1.100000 11.750000 929.200000 12.650000 ;
      RECT 0.000000 10.210000 929.200000 11.750000 ;
      RECT 0.000000 9.310000 928.100000 10.210000 ;
      RECT 0.000000 8.990000 929.200000 9.310000 ;
      RECT 1.100000 8.090000 929.200000 8.990000 ;
      RECT 0.000000 1.100000 929.200000 8.090000 ;
      RECT 1.140000 0.000000 929.200000 1.100000 ;
      RECT 0.000000 0.000000 0.240000 1.100000 ;
    LAYER met4 ;
      RECT 0.000000 918.920000 929.200000 920.720000 ;
      RECT 4.360000 914.920000 924.840000 918.920000 ;
      RECT 923.440000 5.800000 924.840000 914.920000 ;
      RECT 8.360000 5.800000 920.840000 914.920000 ;
      RECT 4.360000 5.800000 5.760000 914.920000 ;
      RECT 927.440000 1.800000 929.200000 918.920000 ;
      RECT 4.360000 1.800000 924.840000 5.800000 ;
      RECT 0.000000 1.800000 1.760000 918.920000 ;
      RECT 0.000000 0.000000 929.200000 1.800000 ;
  END
END user_proj_example

END LIBRARY
