##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Sat Jun 25 21:49:29 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_proj_example
  CLASS BLOCK ;
  SIZE 926.440000 BY 923.440000 ;
  FOREIGN user_proj_example 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9555 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.852 LAYER met4  ;
    ANTENNAMAXAREACAR 4.65704 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 27.0481 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.154225 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1.825000 0.000000 1.965000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3339 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 80.3208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 428.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.455 LAYER met4  ;
    ANTENNAMAXAREACAR 22.3755 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 116.846 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.121796 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1.080000 0.000000 1.220000 0.490000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.905000 0.000000 197.045000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.220000 0.000000 66.360000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.800000 0.000000 198.940000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.010000 0.000000 195.150000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.120000 0.000000 193.260000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.225000 0.000000 191.365000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.330000 0.000000 189.470000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.830000 0.000000 126.970000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.935000 0.000000 125.075000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.040000 0.000000 123.180000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.145000 0.000000 121.285000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.250000 0.000000 119.390000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.360000 0.000000 117.500000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.465000 0.000000 115.605000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.570000 0.000000 113.710000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.675000 0.000000 111.815000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.780000 0.000000 109.920000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.890000 0.000000 108.030000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.995000 0.000000 106.135000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.100000 0.000000 104.240000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.205000 0.000000 102.345000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.310000 0.000000 100.450000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.420000 0.000000 98.560000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.525000 0.000000 96.665000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.630000 0.000000 94.770000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.735000 0.000000 92.875000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.840000 0.000000 90.980000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.950000 0.000000 89.090000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.055000 0.000000 87.195000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.160000 0.000000 85.300000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.265000 0.000000 83.405000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.370000 0.000000 81.510000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.480000 0.000000 79.620000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.585000 0.000000 77.725000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.690000 0.000000 75.830000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.795000 0.000000 73.935000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.900000 0.000000 72.040000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010000 0.000000 70.150000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.115000 0.000000 68.255000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.325000 0.000000 64.465000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.430000 0.000000 62.570000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.540000 0.000000 60.680000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.645000 0.000000 58.785000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.750000 0.000000 56.890000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.855000 0.000000 54.995000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.960000 0.000000 53.100000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.070000 0.000000 51.210000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.175000 0.000000 49.315000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.280000 0.000000 47.420000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.385000 0.000000 45.525000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.490000 0.000000 43.630000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.600000 0.000000 41.740000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.705000 0.000000 39.845000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810000 0.000000 37.950000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.915000 0.000000 36.055000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.020000 0.000000 34.160000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.130000 0.000000 32.270000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.235000 0.000000 30.375000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.340000 0.000000 28.480000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.445000 0.000000 26.585000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.550000 0.000000 24.690000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.660000 0.000000 22.800000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.765000 0.000000 20.905000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.870000 0.000000 19.010000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.975000 0.000000 17.115000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.080000 0.000000 15.220000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.190000 0.000000 13.330000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.295000 0.000000 11.435000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.400000 0.000000 9.540000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.505000 0.000000 7.645000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610000 0.000000 5.750000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2639 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 3.720000 0.000000 3.860000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.8084 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.66 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 187.435000 0.000000 187.575000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 185.540000 0.000000 185.680000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 183.650000 0.000000 183.790000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 181.755000 0.000000 181.895000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 179.860000 0.000000 180.000000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 177.965000 0.000000 178.105000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 176.070000 0.000000 176.210000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 174.180000 0.000000 174.320000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 172.285000 0.000000 172.425000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 170.390000 0.000000 170.530000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 168.495000 0.000000 168.635000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 166.600000 0.000000 166.740000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 164.710000 0.000000 164.850000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 162.815000 0.000000 162.955000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 160.920000 0.000000 161.060000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 159.025000 0.000000 159.165000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 157.130000 0.000000 157.270000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 155.240000 0.000000 155.380000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 153.345000 0.000000 153.485000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 151.450000 0.000000 151.590000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 149.555000 0.000000 149.695000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 147.660000 0.000000 147.800000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 145.770000 0.000000 145.910000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 143.875000 0.000000 144.015000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 141.980000 0.000000 142.120000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 140.085000 0.000000 140.225000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 138.190000 0.000000 138.330000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 136.300000 0.000000 136.440000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 134.405000 0.000000 134.545000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 132.510000 0.000000 132.650000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 130.615000 0.000000 130.755000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 128.720000 0.000000 128.860000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230000 0.000000 441.370000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.340000 0.000000 439.480000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.445000 0.000000 437.585000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.550000 0.000000 435.690000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.655000 0.000000 433.795000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.760000 0.000000 431.900000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.870000 0.000000 430.010000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.975000 0.000000 428.115000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.080000 0.000000 426.220000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.185000 0.000000 424.325000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.290000 0.000000 422.430000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.400000 0.000000 420.540000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.505000 0.000000 418.645000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.610000 0.000000 416.750000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.715000 0.000000 414.855000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.820000 0.000000 412.960000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.930000 0.000000 411.070000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.035000 0.000000 409.175000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.140000 0.000000 407.280000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.245000 0.000000 405.385000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.350000 0.000000 403.490000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.460000 0.000000 401.600000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.565000 0.000000 399.705000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.670000 0.000000 397.810000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.775000 0.000000 395.915000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.880000 0.000000 394.020000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.990000 0.000000 392.130000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.095000 0.000000 390.235000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.200000 0.000000 388.340000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.305000 0.000000 386.445000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.410000 0.000000 384.550000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.520000 0.000000 382.660000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.625000 0.000000 380.765000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.730000 0.000000 378.870000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.835000 0.000000 376.975000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.940000 0.000000 375.080000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.050000 0.000000 373.190000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.155000 0.000000 371.295000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.260000 0.000000 369.400000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.365000 0.000000 367.505000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.470000 0.000000 365.610000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.580000 0.000000 363.720000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.685000 0.000000 361.825000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.790000 0.000000 359.930000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.895000 0.000000 358.035000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.000000 0.000000 356.140000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.110000 0.000000 354.250000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.215000 0.000000 352.355000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.320000 0.000000 350.460000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.425000 0.000000 348.565000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.530000 0.000000 346.670000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.640000 0.000000 344.780000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.745000 0.000000 342.885000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.850000 0.000000 340.990000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.955000 0.000000 339.095000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.060000 0.000000 337.200000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.170000 0.000000 335.310000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.275000 0.000000 333.415000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.380000 0.000000 331.520000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.485000 0.000000 329.625000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.590000 0.000000 327.730000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.700000 0.000000 325.840000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.246 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.299 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 113.633 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 611.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 21.0375 LAYER met4  ;
    ANTENNAMAXAREACAR 68.5875 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 364.187 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 323.805000 0.000000 323.945000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 340.881 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1824.59 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 14.5155 LAYER met4  ;
    ANTENNAMAXAREACAR 104.168 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 532.514 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 321.910000 0.000000 322.050000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.015000 0.000000 320.155000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.120000 0.000000 318.260000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.230000 0.000000 316.370000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.335000 0.000000 314.475000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.440000 0.000000 312.580000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.545000 0.000000 310.685000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.650000 0.000000 308.790000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.760000 0.000000 306.900000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.865000 0.000000 305.005000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.970000 0.000000 303.110000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.075000 0.000000 301.215000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.180000 0.000000 299.320000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.290000 0.000000 297.430000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.395000 0.000000 295.535000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.500000 0.000000 293.640000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.605000 0.000000 291.745000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.710000 0.000000 289.850000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.820000 0.000000 287.960000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.925000 0.000000 286.065000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.030000 0.000000 284.170000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.135000 0.000000 282.275000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.240000 0.000000 280.380000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.350000 0.000000 278.490000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.455000 0.000000 276.595000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.560000 0.000000 274.700000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.665000 0.000000 272.805000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.770000 0.000000 270.910000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.880000 0.000000 269.020000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.985000 0.000000 267.125000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.090000 0.000000 265.230000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.195000 0.000000 263.335000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.300000 0.000000 261.440000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.542 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 14.9876 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.4895 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 259.410000 0.000000 259.550000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0665 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 8.05525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.7934 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.149293 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 257.515000 0.000000 257.655000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.141 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.63872 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.6519 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.147071 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 255.620000 0.000000 255.760000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.801 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 12.6744 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 55.1207 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 253.725000 0.000000 253.865000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7645 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 7.5922 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.1734 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 251.830000 0.000000 251.970000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2745 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 10.3398 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.3274 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 249.940000 0.000000 250.080000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7753 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 6.9703 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.5687 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 248.045000 0.000000 248.185000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.297 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 5.38897 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.137 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 246.150000 0.000000 246.290000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.595 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 7.78869 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.4687 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 244.255000 0.000000 244.395000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2555 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1595 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 11.2559 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.9516 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 242.360000 0.000000 242.500000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.387 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 6.15546 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.9178 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.144803 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 240.470000 0.000000 240.610000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.048 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.05253 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.6579 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 238.575000 0.000000 238.715000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.64 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.092 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 2.69442 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.9293 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.134949 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 236.680000 0.000000 236.820000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1927 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6295 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 5.16346 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.8033 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 234.785000 0.000000 234.925000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.001 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 10.6776 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.899 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 232.890000 0.000000 233.030000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1048 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.19 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.65589 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.7973 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 231.000000 0.000000 231.140000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.105000 0.000000 229.245000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.210000 0.000000 227.350000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.315000 0.000000 225.455000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.420000 0.000000 223.560000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.530000 0.000000 221.670000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.635000 0.000000 219.775000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.740000 0.000000 217.880000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.845000 0.000000 215.985000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.950000 0.000000 214.090000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.060000 0.000000 212.200000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.165000 0.000000 210.305000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.270000 0.000000 208.410000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.375000 0.000000 206.515000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.480000 0.000000 204.620000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.135 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 20.3264 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 98.3818 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 202.590000 0.000000 202.730000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.695000 0.000000 200.835000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.001 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 132.115 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 655.282 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.241315 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 683.665000 0.000000 683.805000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 681.770000 0.000000 681.910000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 679.875000 0.000000 680.015000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 677.980000 0.000000 678.120000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 676.090000 0.000000 676.230000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 674.195000 0.000000 674.335000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 672.300000 0.000000 672.440000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 670.405000 0.000000 670.545000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 668.510000 0.000000 668.650000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 666.620000 0.000000 666.760000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 664.725000 0.000000 664.865000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 662.830000 0.000000 662.970000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 660.935000 0.000000 661.075000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 659.040000 0.000000 659.180000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 657.150000 0.000000 657.290000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 655.255000 0.000000 655.395000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 653.360000 0.000000 653.500000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 651.465000 0.000000 651.605000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 649.570000 0.000000 649.710000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 647.680000 0.000000 647.820000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 645.785000 0.000000 645.925000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 643.890000 0.000000 644.030000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 641.995000 0.000000 642.135000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 640.100000 0.000000 640.240000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 638.210000 0.000000 638.350000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 636.315000 0.000000 636.455000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 634.420000 0.000000 634.560000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 632.525000 0.000000 632.665000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 630.630000 0.000000 630.770000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 628.740000 0.000000 628.880000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 626.845000 0.000000 626.985000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 624.950000 0.000000 625.090000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 623.055000 0.000000 623.195000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 621.160000 0.000000 621.300000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 619.270000 0.000000 619.410000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 617.375000 0.000000 617.515000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 615.480000 0.000000 615.620000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 613.585000 0.000000 613.725000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 611.690000 0.000000 611.830000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 609.800000 0.000000 609.940000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 607.905000 0.000000 608.045000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 606.010000 0.000000 606.150000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 604.115000 0.000000 604.255000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 602.220000 0.000000 602.360000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 600.330000 0.000000 600.470000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 598.435000 0.000000 598.575000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 596.540000 0.000000 596.680000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 594.645000 0.000000 594.785000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 592.750000 0.000000 592.890000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 590.860000 0.000000 591.000000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 588.965000 0.000000 589.105000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 587.070000 0.000000 587.210000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 585.175000 0.000000 585.315000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 583.280000 0.000000 583.420000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 581.390000 0.000000 581.530000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 579.495000 0.000000 579.635000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 577.600000 0.000000 577.740000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 575.705000 0.000000 575.845000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 573.810000 0.000000 573.950000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 571.920000 0.000000 572.060000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 570.025000 0.000000 570.165000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 568.130000 0.000000 568.270000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.102 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.671 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 566.235000 0.000000 566.375000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.001 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.861 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 564.340000 0.000000 564.480000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.431 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 98.6538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 526.624 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 562.450000 0.000000 562.590000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 85.6128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 457.072 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 560.555000 0.000000 560.695000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 85.7238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 457.664 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 558.660000 0.000000 558.800000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3639 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.58 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 91.3566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.176 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 556.765000 0.000000 556.905000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.752 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 75.6186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 404.24 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 554.870000 0.000000 555.010000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.721 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.0776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 502.688 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 552.980000 0.000000 553.120000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7598 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.638 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.817 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 83.0268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 443.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 551.085000 0.000000 551.225000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.616 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 75.9528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 405.552 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 549.190000 0.000000 549.330000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5564 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.621 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.092 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 83.1228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 443.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 547.295000 0.000000 547.435000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5512 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 96.5688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 515.504 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 545.400000 0.000000 545.540000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5442 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.56 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.071 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 82.4538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 440.224 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 543.510000 0.000000 543.650000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.862 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.101 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 72.3018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 386.08 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 541.615000 0.000000 541.755000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 99.6168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 531.76 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 539.720000 0.000000 539.860000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.192 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.241 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 84.8328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 452.912 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 537.825000 0.000000 537.965000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8467 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.0725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.792 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 72.3408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 386.288 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 535.930000 0.000000 536.070000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.9395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 87.7368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 468.4 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 534.040000 0.000000 534.180000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.68 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 92.7966 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 495.856 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 532.145000 0.000000 532.285000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3921 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.7995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 89.5758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 478.208 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 530.250000 0.000000 530.390000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6668 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.173 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 71.6328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 382.512 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 528.355000 0.000000 528.495000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9385 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 101.693 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 542.832 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 526.460000 0.000000 526.600000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7185 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.238 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 104.9 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 559.936 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 524.570000 0.000000 524.710000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9652 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.547 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 87.4188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 466.704 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 522.675000 0.000000 522.815000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.47 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 99.6798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 532.096 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 520.780000 0.000000 520.920000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3611 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.344 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.515 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 99.5754 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 532.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 518.885000 0.000000 519.025000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.1605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.137 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 96.9906 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 518.224 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 516.990000 0.000000 517.130000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 100.412 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 536 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 515.100000 0.000000 515.240000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.416 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.4746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 419.472 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 513.205000 0.000000 513.345000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6233 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.653 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 101.947 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 544.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 511.310000 0.000000 511.450000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 100.468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 536.768 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 509.415000 0.000000 509.555000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5932 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.7466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 506.256 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 507.520000 0.000000 507.660000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9077 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 100.826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 538.208 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 505.630000 0.000000 505.770000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.513 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.389 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 100.85 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 538.336 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 503.735000 0.000000 503.875000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.001 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.861 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 501.840000 0.000000 501.980000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 499.945000 0.000000 500.085000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 498.050000 0.000000 498.190000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 496.160000 0.000000 496.300000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.4767 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.172 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 128.999 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 494.265000 0.000000 494.405000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.779 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.488 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 492.370000 0.000000 492.510000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 490.475000 0.000000 490.615000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 488.580000 0.000000 488.720000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 486.690000 0.000000 486.830000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 484.795000 0.000000 484.935000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 482.900000 0.000000 483.040000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 481.005000 0.000000 481.145000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 479.110000 0.000000 479.250000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 477.220000 0.000000 477.360000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 475.325000 0.000000 475.465000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 473.430000 0.000000 473.570000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 471.535000 0.000000 471.675000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 469.640000 0.000000 469.780000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 467.750000 0.000000 467.890000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 465.855000 0.000000 465.995000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 463.960000 0.000000 464.100000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 462.065000 0.000000 462.205000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 460.170000 0.000000 460.310000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 458.280000 0.000000 458.420000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 456.385000 0.000000 456.525000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 454.490000 0.000000 454.630000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 452.595000 0.000000 452.735000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 450.700000 0.000000 450.840000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 448.810000 0.000000 448.950000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.537 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 446.915000 0.000000 447.055000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.7888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 445.020000 0.000000 445.160000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.8084 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.66 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 443.125000 0.000000 443.265000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.095000 0.000000 926.235000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.200000 0.000000 924.340000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.310000 0.000000 922.450000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.415000 0.000000 920.555000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.520000 0.000000 918.660000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.625000 0.000000 916.765000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.730000 0.000000 914.870000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.840000 0.000000 912.980000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.945000 0.000000 911.085000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.050000 0.000000 909.190000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.155000 0.000000 907.295000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.260000 0.000000 905.400000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.370000 0.000000 903.510000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.475000 0.000000 901.615000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.580000 0.000000 899.720000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.685000 0.000000 897.825000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.790000 0.000000 895.930000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.900000 0.000000 894.040000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.005000 0.000000 892.145000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.110000 0.000000 890.250000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.215000 0.000000 888.355000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.320000 0.000000 886.460000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.430000 0.000000 884.570000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.535000 0.000000 882.675000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.640000 0.000000 880.780000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.745000 0.000000 878.885000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.850000 0.000000 876.990000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.960000 0.000000 875.100000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.065000 0.000000 873.205000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.170000 0.000000 871.310000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.275000 0.000000 869.415000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.380000 0.000000 867.520000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.490000 0.000000 865.630000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.595000 0.000000 863.735000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.700000 0.000000 861.840000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.805000 0.000000 859.945000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.910000 0.000000 858.050000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.020000 0.000000 856.160000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.125000 0.000000 854.265000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.230000 0.000000 852.370000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.335000 0.000000 850.475000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.440000 0.000000 848.580000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.550000 0.000000 846.690000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.655000 0.000000 844.795000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.760000 0.000000 842.900000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.865000 0.000000 841.005000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.970000 0.000000 839.110000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.080000 0.000000 837.220000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.185000 0.000000 835.325000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.290000 0.000000 833.430000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.395000 0.000000 831.535000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.500000 0.000000 829.640000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.610000 0.000000 827.750000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.715000 0.000000 825.855000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.820000 0.000000 823.960000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.925000 0.000000 822.065000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.030000 0.000000 820.170000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.140000 0.000000 818.280000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.245000 0.000000 816.385000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.350000 0.000000 814.490000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.455000 0.000000 812.595000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.560000 0.000000 810.700000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 288.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 124.283 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 668 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 34.308 LAYER met4  ;
    ANTENNAMAXAREACAR 12.9056 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 66.8518 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.132727 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 808.670000 0.000000 808.810000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.655 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.114 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.54 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 650.799 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3478.9 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 21.9405 LAYER met4  ;
    ANTENNAMAXAREACAR 65.5369 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 345.459 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.289249 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 806.775000 0.000000 806.915000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.714 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 15.877 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.4325 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 804.880000 0.000000 805.020000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6205 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.5012 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.254 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 802.985000 0.000000 803.125000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.575 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.9873 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.9325 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 801.090000 0.000000 801.230000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.696 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.372 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 20.0444 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.9564 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 799.200000 0.000000 799.340000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9065 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.623 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.627 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 797.305000 0.000000 797.445000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.323 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.4472 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.4484 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 795.410000 0.000000 795.550000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5225 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 16.9746 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.4048 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 793.515000 0.000000 793.655000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6624 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.204 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.2222 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.8452 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 791.620000 0.000000 791.760000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5686 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.735 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 20.3952 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.4881 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 789.730000 0.000000 789.870000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1725 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 20.2528 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.4762 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 787.835000 0.000000 787.975000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.696 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.372 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.6651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.3214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 785.940000 0.000000 786.080000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4175 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 16.654 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.5397 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 784.045000 0.000000 784.185000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.924 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.1397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.2103 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 782.150000 0.000000 782.290000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.344 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.9694 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.0595 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 780.260000 0.000000 780.400000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1445 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 16.3746 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.4048 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 778.365000 0.000000 778.505000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7058 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.421 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.0778 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.123 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 776.470000 0.000000 776.610000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5721 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7525 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.8675 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.8492 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 774.575000 0.000000 774.715000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.19 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.725 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.8373 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 772.680000 0.000000 772.820000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.295 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 16.6135 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.5992 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 770.790000 0.000000 770.930000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5715 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.3167 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.3175 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 768.895000 0.000000 769.035000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.542 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.602 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 15.6992 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.5436 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 767.000000 0.000000 767.140000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0885 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.5639 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.0317 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 765.105000 0.000000 765.245000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.302 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 19.1651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 84.8214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 763.210000 0.000000 763.350000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7492 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.638 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 20.9778 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 94.623 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 761.320000 0.000000 761.460000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5763 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7735 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.3897 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.4603 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 759.425000 0.000000 759.565000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6638 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.211 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.2472 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.4484 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 757.530000 0.000000 757.670000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.366 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.3135 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.0992 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 755.635000 0.000000 755.775000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7324 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.554 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.7341 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 753.740000 0.000000 753.880000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.623 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 15.7325 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.7103 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 751.850000 0.000000 751.990000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 19.575 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.0873 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 749.955000 0.000000 750.095000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.344 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 22.1984 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 99.9881 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 748.060000 0.000000 748.200000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6205 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 25.0389 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 114.929 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 746.165000 0.000000 746.305000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.183 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.12343 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.6434 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 744.270000 0.000000 744.410000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.018 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.982 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.7503 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.9162 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 742.380000 0.000000 742.520000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7247 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5155 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 3.89677 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.6465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 740.485000 0.000000 740.625000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4142 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.963 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 5.3905 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.9788 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 738.590000 0.000000 738.730000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1165 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 3.73556 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.8404 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 736.695000 0.000000 736.835000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9704 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.744 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.88424 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.4475 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 734.800000 0.000000 734.940000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6946 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.365 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 3.83596 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.3424 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 732.910000 0.000000 733.050000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3475 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.1899 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.9758 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 731.015000 0.000000 731.155000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6792 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.16586 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.8556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 729.120000 0.000000 729.260000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2495 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.0202 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.1273 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 727.225000 0.000000 727.365000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.877 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.44687 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.397 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 725.330000 0.000000 725.470000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9676 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.73 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.79374 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.9949 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 723.440000 0.000000 723.580000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6225 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 5.54545 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.7556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 721.545000 0.000000 721.685000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6414 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.099 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 3.72848 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.805 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 719.650000 0.000000 719.790000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8935 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.09717 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.4101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 717.755000 0.000000 717.895000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.01 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.86162 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.3343 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 715.860000 0.000000 716.000000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.970000 0.000000 714.110000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.075000 0.000000 712.215000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.180000 0.000000 710.320000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.285000 0.000000 708.425000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.390000 0.000000 706.530000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.500000 0.000000 704.640000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.605000 0.000000 702.745000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.710000 0.000000 700.850000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.815000 0.000000 698.955000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.920000 0.000000 697.060000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.030000 0.000000 695.170000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.135000 0.000000 693.275000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.240000 0.000000 691.380000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.345000 0.000000 689.485000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.866 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 11.8414 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.4051 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 687.450000 0.000000 687.590000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.560000 0.000000 685.700000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 44.895000 0.800000 45.195000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 112.460000 0.800000 112.760000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 180.025000 0.800000 180.325000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 247.590000 0.800000 247.890000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 315.160000 0.800000 315.460000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 382.725000 0.800000 383.025000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 450.290000 0.800000 450.590000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 517.855000 0.800000 518.155000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 585.420000 0.800000 585.720000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 652.990000 0.800000 653.290000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 720.555000 0.800000 720.855000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 788.120000 0.800000 788.420000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 855.685000 0.800000 855.985000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 919.730000 0.800000 920.030000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.195000 922.950000 71.335000 923.440000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.090000 922.950000 178.230000 923.440000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.985000 922.950000 285.125000 923.440000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.880000 922.950000 392.020000 923.440000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.780000 922.950000 498.920000 923.440000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.675000 922.950000 605.815000 923.440000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.570000 922.950000 712.710000 923.440000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.465000 922.950000 819.605000 923.440000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.480000 922.950000 916.620000 923.440000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 881.305000 926.440000 881.605000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 818.345000 926.440000 818.645000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 755.380000 926.440000 755.680000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 692.420000 926.440000 692.720000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 629.460000 926.440000 629.760000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 566.500000 926.440000 566.800000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 503.540000 926.440000 503.840000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 440.575000 926.440000 440.875000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 377.615000 926.440000 377.915000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2039 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 30.0945 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 154.772 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 314.655000 926.440000 314.955000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 251.695000 926.440000 251.995000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 188.735000 926.440000 189.035000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 125.770000 926.440000 126.070000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 62.810000 926.440000 63.110000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 925.640000 4.730000 926.440000 5.030000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 22.370000 0.800000 22.670000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 129.153 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 689.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 84.8088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 452.784 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 89.940000 0.800000 90.240000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 128.153 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 683.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 83.3448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 444.976 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 157.505000 0.800000 157.805000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 128.097 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 683.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 80.9658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 432.288 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 225.070000 0.800000 225.370000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 114.425 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 610.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.3538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.024 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 292.635000 0.800000 292.935000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 124.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.5326 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.448 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 360.200000 0.800000 360.500000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 126.618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 677.648 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 427.770000 0.800000 428.070000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1891 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 139.293 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 745.248 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 495.335000 0.800000 495.635000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2826 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 286.157 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1527.58 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 562.900000 0.800000 563.200000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9841 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 297.361 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1586.86 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 630.465000 0.800000 630.765000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8116 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 190.915 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1020.1 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 698.030000 0.800000 698.330000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7826 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 330.34 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1762.75 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 765.600000 0.800000 765.900000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.1169 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 108.329 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 578.224 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 833.165000 0.800000 833.465000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8234 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 102.974 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 549.664 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 900.730000 0.800000 901.030000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.3323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 176.382 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 108.815 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 580.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 35.560000 922.950000 35.700000 923.440000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.3537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.6075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.762 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 185.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 231.796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1238.13 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 142.460000 922.950000 142.600000 923.440000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.2 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.437 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 263.641 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1407.97 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 249.355000 922.950000 249.495000 923.440000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.2677 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.1775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 229.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 353.419 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1885.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 356.250000 922.950000 356.390000 923.440000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.0195 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.8715 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 463.145000 922.950000 463.285000 923.440000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 115.351 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 615.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.9718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 160.32 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 570.040000 922.950000 570.180000 923.440000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.0765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.6176 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 201.568 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 676.940000 922.950000 677.080000 923.440000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6515 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 88.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 471.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.0438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 160.704 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 783.835000 922.950000 783.975000 923.440000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6851 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 84.43 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 450.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.5168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 890.730000 922.950000 890.870000 923.440000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.2308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 204.368 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 902.290000 926.440000 902.590000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 83.0974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 443.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.4306 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 189.904 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 839.330000 926.440000 839.630000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 123.259 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 658.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 776.370000 926.440000 776.670000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8054 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.2114 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.872 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 713.410000 926.440000 713.710000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3751 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 81.8712 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 438.528 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 650.445000 926.440000 650.745000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.8002 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 304.816 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 587.485000 926.440000 587.785000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4691 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.5022 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.56 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 524.525000 926.440000 524.825000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2281 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.9316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 160.576 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 461.565000 926.440000 461.865000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 89.2099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 476.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.5628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.472 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 398.605000 926.440000 398.905000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 335.640000 926.440000 335.940000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 78.0316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 416.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.8926 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.368 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 272.680000 926.440000 272.980000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 209.720000 926.440000 210.020000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 146.760000 926.440000 147.060000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5236 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 83.800000 926.440000 84.100000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 67.1897 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 358.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.267017 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 20.835000 926.440000 21.135000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.8399 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.540000 0.000000 0.840000 0.800000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 67.415000 0.800000 67.715000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 134.980000 0.800000 135.280000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 202.550000 0.800000 202.850000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8731 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 270.115000 0.800000 270.415000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 337.680000 0.800000 337.980000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9391 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 405.245000 0.800000 405.545000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9256 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 472.810000 0.800000 473.110000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 540.380000 0.800000 540.680000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8851 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 607.945000 0.800000 608.245000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 675.510000 0.800000 675.810000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met3  ;
    ANTENNAMAXAREACAR 16.2373 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 91.8251 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 139.482 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 751.237 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 743.075000 0.800000 743.375000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met3  ;
    ANTENNAMAXAREACAR 16.2373 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 91.8251 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 139.482 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 751.237 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 810.640000 0.800000 810.940000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met3  ;
    ANTENNAMAXAREACAR 89.6567 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 444.339 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.307193 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 212.901 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1103.75 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.307193 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 878.210000 0.800000 878.510000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4986 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.282 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met3  ;
    ANTENNAMAXAREACAR 16.5463 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 93.4727 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 139.791 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 752.885 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 15.340000 922.950000 15.480000 923.440000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4741 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.1595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met3  ;
    ANTENNAMAXAREACAR 16.5463 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 93.4727 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 139.791 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 752.885 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 106.825000 922.950000 106.965000 923.440000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4741 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.1595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met3  ;
    ANTENNAMAXAREACAR 16.5463 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 93.4727 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 139.791 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 752.885 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 213.720000 922.950000 213.860000 923.440000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4741 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.1595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met3  ;
    ANTENNAMAXAREACAR 16.5463 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 93.4727 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 139.791 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 752.885 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 320.620000 922.950000 320.760000 923.440000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.0125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met3  ;
    ANTENNAMAXAREACAR 16.5463 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 93.4727 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 139.791 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 752.885 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0633714 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 427.515000 922.950000 427.655000 923.440000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 56.1479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 279.562 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.28 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.8849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 534.410000 922.950000 534.550000 923.440000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 56.1479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 279.562 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.28 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.8849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 641.305000 922.950000 641.445000 923.440000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 56.1479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 279.562 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.28 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.8849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 748.200000 922.950000 748.340000 923.440000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 56.1381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 279.415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.28 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.8849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 855.100000 922.950000 855.240000 923.440000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7649 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 919.730000 926.440000 920.030000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6899 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 860.315000 926.440000 860.615000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7649 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 797.355000 926.440000 797.655000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6899 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 734.395000 926.440000 734.695000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6899 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 671.435000 926.440000 671.735000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6899 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 608.475000 926.440000 608.775000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6449 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 545.510000 926.440000 545.810000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 482.550000 926.440000 482.850000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 419.590000 926.440000 419.890000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.744 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 356.630000 926.440000 356.930000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 293.670000 926.440000 293.970000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2941 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 230.705000 926.440000 231.005000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4531 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 167.745000 926.440000 168.045000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2161 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 104.785000 926.440000 105.085000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3601 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 161.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 866.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3134 LAYER met4  ;
    ANTENNAMAXAREACAR 123.244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.412 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 925.640000 41.825000 926.440000 42.125000 ;
    END
  END io_oeb[0]
  PIN irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 15.100000 0.800000 15.400000 ;
    END
  END irq[2]
  PIN irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 10.220000 0.800000 10.520000 ;
    END
  END irq[1]
  PIN irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 187.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 999.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 5.340000 0.800000 5.640000 ;
    END
  END irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 922.380000 2.100000 924.380000 921.340000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.060000 2.100000 4.060000 921.340000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 434.900000 514.330000 436.640000 909.110000 ;
      LAYER met4 ;
        RECT 910.220000 514.330000 911.960000 909.110000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 918.380000 6.100000 920.380000 917.340000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.060000 6.100000 8.060000 917.340000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 906.820000 517.730000 908.560000 905.710000 ;
      LAYER met4 ;
        RECT 438.300000 517.730000 440.040000 905.710000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 926.440000 923.440000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 926.440000 923.440000 ;
    LAYER met2 ;
      RECT 916.760000 922.810000 926.440000 923.440000 ;
      RECT 891.010000 922.810000 916.340000 923.440000 ;
      RECT 855.380000 922.810000 890.590000 923.440000 ;
      RECT 819.745000 922.810000 854.960000 923.440000 ;
      RECT 784.115000 922.810000 819.325000 923.440000 ;
      RECT 748.480000 922.810000 783.695000 923.440000 ;
      RECT 712.850000 922.810000 748.060000 923.440000 ;
      RECT 677.220000 922.810000 712.430000 923.440000 ;
      RECT 641.585000 922.810000 676.800000 923.440000 ;
      RECT 605.955000 922.810000 641.165000 923.440000 ;
      RECT 570.320000 922.810000 605.535000 923.440000 ;
      RECT 534.690000 922.810000 569.900000 923.440000 ;
      RECT 499.060000 922.810000 534.270000 923.440000 ;
      RECT 463.425000 922.810000 498.640000 923.440000 ;
      RECT 427.795000 922.810000 463.005000 923.440000 ;
      RECT 392.160000 922.810000 427.375000 923.440000 ;
      RECT 356.530000 922.810000 391.740000 923.440000 ;
      RECT 320.900000 922.810000 356.110000 923.440000 ;
      RECT 285.265000 922.810000 320.480000 923.440000 ;
      RECT 249.635000 922.810000 284.845000 923.440000 ;
      RECT 214.000000 922.810000 249.215000 923.440000 ;
      RECT 178.370000 922.810000 213.580000 923.440000 ;
      RECT 142.740000 922.810000 177.950000 923.440000 ;
      RECT 107.105000 922.810000 142.320000 923.440000 ;
      RECT 71.475000 922.810000 106.685000 923.440000 ;
      RECT 35.840000 922.810000 71.055000 923.440000 ;
      RECT 15.620000 922.810000 35.420000 923.440000 ;
      RECT 0.000000 922.810000 15.200000 923.440000 ;
      RECT 0.000000 0.630000 926.440000 922.810000 ;
      RECT 926.375000 0.000000 926.440000 0.630000 ;
      RECT 924.480000 0.000000 925.955000 0.630000 ;
      RECT 922.590000 0.000000 924.060000 0.630000 ;
      RECT 920.695000 0.000000 922.170000 0.630000 ;
      RECT 918.800000 0.000000 920.275000 0.630000 ;
      RECT 916.905000 0.000000 918.380000 0.630000 ;
      RECT 915.010000 0.000000 916.485000 0.630000 ;
      RECT 913.120000 0.000000 914.590000 0.630000 ;
      RECT 911.225000 0.000000 912.700000 0.630000 ;
      RECT 909.330000 0.000000 910.805000 0.630000 ;
      RECT 907.435000 0.000000 908.910000 0.630000 ;
      RECT 905.540000 0.000000 907.015000 0.630000 ;
      RECT 903.650000 0.000000 905.120000 0.630000 ;
      RECT 901.755000 0.000000 903.230000 0.630000 ;
      RECT 899.860000 0.000000 901.335000 0.630000 ;
      RECT 897.965000 0.000000 899.440000 0.630000 ;
      RECT 896.070000 0.000000 897.545000 0.630000 ;
      RECT 894.180000 0.000000 895.650000 0.630000 ;
      RECT 892.285000 0.000000 893.760000 0.630000 ;
      RECT 890.390000 0.000000 891.865000 0.630000 ;
      RECT 888.495000 0.000000 889.970000 0.630000 ;
      RECT 886.600000 0.000000 888.075000 0.630000 ;
      RECT 884.710000 0.000000 886.180000 0.630000 ;
      RECT 882.815000 0.000000 884.290000 0.630000 ;
      RECT 880.920000 0.000000 882.395000 0.630000 ;
      RECT 879.025000 0.000000 880.500000 0.630000 ;
      RECT 877.130000 0.000000 878.605000 0.630000 ;
      RECT 875.240000 0.000000 876.710000 0.630000 ;
      RECT 873.345000 0.000000 874.820000 0.630000 ;
      RECT 871.450000 0.000000 872.925000 0.630000 ;
      RECT 869.555000 0.000000 871.030000 0.630000 ;
      RECT 867.660000 0.000000 869.135000 0.630000 ;
      RECT 865.770000 0.000000 867.240000 0.630000 ;
      RECT 863.875000 0.000000 865.350000 0.630000 ;
      RECT 861.980000 0.000000 863.455000 0.630000 ;
      RECT 860.085000 0.000000 861.560000 0.630000 ;
      RECT 858.190000 0.000000 859.665000 0.630000 ;
      RECT 856.300000 0.000000 857.770000 0.630000 ;
      RECT 854.405000 0.000000 855.880000 0.630000 ;
      RECT 852.510000 0.000000 853.985000 0.630000 ;
      RECT 850.615000 0.000000 852.090000 0.630000 ;
      RECT 848.720000 0.000000 850.195000 0.630000 ;
      RECT 846.830000 0.000000 848.300000 0.630000 ;
      RECT 844.935000 0.000000 846.410000 0.630000 ;
      RECT 843.040000 0.000000 844.515000 0.630000 ;
      RECT 841.145000 0.000000 842.620000 0.630000 ;
      RECT 839.250000 0.000000 840.725000 0.630000 ;
      RECT 837.360000 0.000000 838.830000 0.630000 ;
      RECT 835.465000 0.000000 836.940000 0.630000 ;
      RECT 833.570000 0.000000 835.045000 0.630000 ;
      RECT 831.675000 0.000000 833.150000 0.630000 ;
      RECT 829.780000 0.000000 831.255000 0.630000 ;
      RECT 827.890000 0.000000 829.360000 0.630000 ;
      RECT 825.995000 0.000000 827.470000 0.630000 ;
      RECT 824.100000 0.000000 825.575000 0.630000 ;
      RECT 822.205000 0.000000 823.680000 0.630000 ;
      RECT 820.310000 0.000000 821.785000 0.630000 ;
      RECT 818.420000 0.000000 819.890000 0.630000 ;
      RECT 816.525000 0.000000 818.000000 0.630000 ;
      RECT 814.630000 0.000000 816.105000 0.630000 ;
      RECT 812.735000 0.000000 814.210000 0.630000 ;
      RECT 810.840000 0.000000 812.315000 0.630000 ;
      RECT 808.950000 0.000000 810.420000 0.630000 ;
      RECT 807.055000 0.000000 808.530000 0.630000 ;
      RECT 805.160000 0.000000 806.635000 0.630000 ;
      RECT 803.265000 0.000000 804.740000 0.630000 ;
      RECT 801.370000 0.000000 802.845000 0.630000 ;
      RECT 799.480000 0.000000 800.950000 0.630000 ;
      RECT 797.585000 0.000000 799.060000 0.630000 ;
      RECT 795.690000 0.000000 797.165000 0.630000 ;
      RECT 793.795000 0.000000 795.270000 0.630000 ;
      RECT 791.900000 0.000000 793.375000 0.630000 ;
      RECT 790.010000 0.000000 791.480000 0.630000 ;
      RECT 788.115000 0.000000 789.590000 0.630000 ;
      RECT 786.220000 0.000000 787.695000 0.630000 ;
      RECT 784.325000 0.000000 785.800000 0.630000 ;
      RECT 782.430000 0.000000 783.905000 0.630000 ;
      RECT 780.540000 0.000000 782.010000 0.630000 ;
      RECT 778.645000 0.000000 780.120000 0.630000 ;
      RECT 776.750000 0.000000 778.225000 0.630000 ;
      RECT 774.855000 0.000000 776.330000 0.630000 ;
      RECT 772.960000 0.000000 774.435000 0.630000 ;
      RECT 771.070000 0.000000 772.540000 0.630000 ;
      RECT 769.175000 0.000000 770.650000 0.630000 ;
      RECT 767.280000 0.000000 768.755000 0.630000 ;
      RECT 765.385000 0.000000 766.860000 0.630000 ;
      RECT 763.490000 0.000000 764.965000 0.630000 ;
      RECT 761.600000 0.000000 763.070000 0.630000 ;
      RECT 759.705000 0.000000 761.180000 0.630000 ;
      RECT 757.810000 0.000000 759.285000 0.630000 ;
      RECT 755.915000 0.000000 757.390000 0.630000 ;
      RECT 754.020000 0.000000 755.495000 0.630000 ;
      RECT 752.130000 0.000000 753.600000 0.630000 ;
      RECT 750.235000 0.000000 751.710000 0.630000 ;
      RECT 748.340000 0.000000 749.815000 0.630000 ;
      RECT 746.445000 0.000000 747.920000 0.630000 ;
      RECT 744.550000 0.000000 746.025000 0.630000 ;
      RECT 742.660000 0.000000 744.130000 0.630000 ;
      RECT 740.765000 0.000000 742.240000 0.630000 ;
      RECT 738.870000 0.000000 740.345000 0.630000 ;
      RECT 736.975000 0.000000 738.450000 0.630000 ;
      RECT 735.080000 0.000000 736.555000 0.630000 ;
      RECT 733.190000 0.000000 734.660000 0.630000 ;
      RECT 731.295000 0.000000 732.770000 0.630000 ;
      RECT 729.400000 0.000000 730.875000 0.630000 ;
      RECT 727.505000 0.000000 728.980000 0.630000 ;
      RECT 725.610000 0.000000 727.085000 0.630000 ;
      RECT 723.720000 0.000000 725.190000 0.630000 ;
      RECT 721.825000 0.000000 723.300000 0.630000 ;
      RECT 719.930000 0.000000 721.405000 0.630000 ;
      RECT 718.035000 0.000000 719.510000 0.630000 ;
      RECT 716.140000 0.000000 717.615000 0.630000 ;
      RECT 714.250000 0.000000 715.720000 0.630000 ;
      RECT 712.355000 0.000000 713.830000 0.630000 ;
      RECT 710.460000 0.000000 711.935000 0.630000 ;
      RECT 708.565000 0.000000 710.040000 0.630000 ;
      RECT 706.670000 0.000000 708.145000 0.630000 ;
      RECT 704.780000 0.000000 706.250000 0.630000 ;
      RECT 702.885000 0.000000 704.360000 0.630000 ;
      RECT 700.990000 0.000000 702.465000 0.630000 ;
      RECT 699.095000 0.000000 700.570000 0.630000 ;
      RECT 697.200000 0.000000 698.675000 0.630000 ;
      RECT 695.310000 0.000000 696.780000 0.630000 ;
      RECT 693.415000 0.000000 694.890000 0.630000 ;
      RECT 691.520000 0.000000 692.995000 0.630000 ;
      RECT 689.625000 0.000000 691.100000 0.630000 ;
      RECT 687.730000 0.000000 689.205000 0.630000 ;
      RECT 685.840000 0.000000 687.310000 0.630000 ;
      RECT 683.945000 0.000000 685.420000 0.630000 ;
      RECT 682.050000 0.000000 683.525000 0.630000 ;
      RECT 680.155000 0.000000 681.630000 0.630000 ;
      RECT 678.260000 0.000000 679.735000 0.630000 ;
      RECT 676.370000 0.000000 677.840000 0.630000 ;
      RECT 674.475000 0.000000 675.950000 0.630000 ;
      RECT 672.580000 0.000000 674.055000 0.630000 ;
      RECT 670.685000 0.000000 672.160000 0.630000 ;
      RECT 668.790000 0.000000 670.265000 0.630000 ;
      RECT 666.900000 0.000000 668.370000 0.630000 ;
      RECT 665.005000 0.000000 666.480000 0.630000 ;
      RECT 663.110000 0.000000 664.585000 0.630000 ;
      RECT 661.215000 0.000000 662.690000 0.630000 ;
      RECT 659.320000 0.000000 660.795000 0.630000 ;
      RECT 657.430000 0.000000 658.900000 0.630000 ;
      RECT 655.535000 0.000000 657.010000 0.630000 ;
      RECT 653.640000 0.000000 655.115000 0.630000 ;
      RECT 651.745000 0.000000 653.220000 0.630000 ;
      RECT 649.850000 0.000000 651.325000 0.630000 ;
      RECT 647.960000 0.000000 649.430000 0.630000 ;
      RECT 646.065000 0.000000 647.540000 0.630000 ;
      RECT 644.170000 0.000000 645.645000 0.630000 ;
      RECT 642.275000 0.000000 643.750000 0.630000 ;
      RECT 640.380000 0.000000 641.855000 0.630000 ;
      RECT 638.490000 0.000000 639.960000 0.630000 ;
      RECT 636.595000 0.000000 638.070000 0.630000 ;
      RECT 634.700000 0.000000 636.175000 0.630000 ;
      RECT 632.805000 0.000000 634.280000 0.630000 ;
      RECT 630.910000 0.000000 632.385000 0.630000 ;
      RECT 629.020000 0.000000 630.490000 0.630000 ;
      RECT 627.125000 0.000000 628.600000 0.630000 ;
      RECT 625.230000 0.000000 626.705000 0.630000 ;
      RECT 623.335000 0.000000 624.810000 0.630000 ;
      RECT 621.440000 0.000000 622.915000 0.630000 ;
      RECT 619.550000 0.000000 621.020000 0.630000 ;
      RECT 617.655000 0.000000 619.130000 0.630000 ;
      RECT 615.760000 0.000000 617.235000 0.630000 ;
      RECT 613.865000 0.000000 615.340000 0.630000 ;
      RECT 611.970000 0.000000 613.445000 0.630000 ;
      RECT 610.080000 0.000000 611.550000 0.630000 ;
      RECT 608.185000 0.000000 609.660000 0.630000 ;
      RECT 606.290000 0.000000 607.765000 0.630000 ;
      RECT 604.395000 0.000000 605.870000 0.630000 ;
      RECT 602.500000 0.000000 603.975000 0.630000 ;
      RECT 600.610000 0.000000 602.080000 0.630000 ;
      RECT 598.715000 0.000000 600.190000 0.630000 ;
      RECT 596.820000 0.000000 598.295000 0.630000 ;
      RECT 594.925000 0.000000 596.400000 0.630000 ;
      RECT 593.030000 0.000000 594.505000 0.630000 ;
      RECT 591.140000 0.000000 592.610000 0.630000 ;
      RECT 589.245000 0.000000 590.720000 0.630000 ;
      RECT 587.350000 0.000000 588.825000 0.630000 ;
      RECT 585.455000 0.000000 586.930000 0.630000 ;
      RECT 583.560000 0.000000 585.035000 0.630000 ;
      RECT 581.670000 0.000000 583.140000 0.630000 ;
      RECT 579.775000 0.000000 581.250000 0.630000 ;
      RECT 577.880000 0.000000 579.355000 0.630000 ;
      RECT 575.985000 0.000000 577.460000 0.630000 ;
      RECT 574.090000 0.000000 575.565000 0.630000 ;
      RECT 572.200000 0.000000 573.670000 0.630000 ;
      RECT 570.305000 0.000000 571.780000 0.630000 ;
      RECT 568.410000 0.000000 569.885000 0.630000 ;
      RECT 566.515000 0.000000 567.990000 0.630000 ;
      RECT 564.620000 0.000000 566.095000 0.630000 ;
      RECT 562.730000 0.000000 564.200000 0.630000 ;
      RECT 560.835000 0.000000 562.310000 0.630000 ;
      RECT 558.940000 0.000000 560.415000 0.630000 ;
      RECT 557.045000 0.000000 558.520000 0.630000 ;
      RECT 555.150000 0.000000 556.625000 0.630000 ;
      RECT 553.260000 0.000000 554.730000 0.630000 ;
      RECT 551.365000 0.000000 552.840000 0.630000 ;
      RECT 549.470000 0.000000 550.945000 0.630000 ;
      RECT 547.575000 0.000000 549.050000 0.630000 ;
      RECT 545.680000 0.000000 547.155000 0.630000 ;
      RECT 543.790000 0.000000 545.260000 0.630000 ;
      RECT 541.895000 0.000000 543.370000 0.630000 ;
      RECT 540.000000 0.000000 541.475000 0.630000 ;
      RECT 538.105000 0.000000 539.580000 0.630000 ;
      RECT 536.210000 0.000000 537.685000 0.630000 ;
      RECT 534.320000 0.000000 535.790000 0.630000 ;
      RECT 532.425000 0.000000 533.900000 0.630000 ;
      RECT 530.530000 0.000000 532.005000 0.630000 ;
      RECT 528.635000 0.000000 530.110000 0.630000 ;
      RECT 526.740000 0.000000 528.215000 0.630000 ;
      RECT 524.850000 0.000000 526.320000 0.630000 ;
      RECT 522.955000 0.000000 524.430000 0.630000 ;
      RECT 521.060000 0.000000 522.535000 0.630000 ;
      RECT 519.165000 0.000000 520.640000 0.630000 ;
      RECT 517.270000 0.000000 518.745000 0.630000 ;
      RECT 515.380000 0.000000 516.850000 0.630000 ;
      RECT 513.485000 0.000000 514.960000 0.630000 ;
      RECT 511.590000 0.000000 513.065000 0.630000 ;
      RECT 509.695000 0.000000 511.170000 0.630000 ;
      RECT 507.800000 0.000000 509.275000 0.630000 ;
      RECT 505.910000 0.000000 507.380000 0.630000 ;
      RECT 504.015000 0.000000 505.490000 0.630000 ;
      RECT 502.120000 0.000000 503.595000 0.630000 ;
      RECT 500.225000 0.000000 501.700000 0.630000 ;
      RECT 498.330000 0.000000 499.805000 0.630000 ;
      RECT 496.440000 0.000000 497.910000 0.630000 ;
      RECT 494.545000 0.000000 496.020000 0.630000 ;
      RECT 492.650000 0.000000 494.125000 0.630000 ;
      RECT 490.755000 0.000000 492.230000 0.630000 ;
      RECT 488.860000 0.000000 490.335000 0.630000 ;
      RECT 486.970000 0.000000 488.440000 0.630000 ;
      RECT 485.075000 0.000000 486.550000 0.630000 ;
      RECT 483.180000 0.000000 484.655000 0.630000 ;
      RECT 481.285000 0.000000 482.760000 0.630000 ;
      RECT 479.390000 0.000000 480.865000 0.630000 ;
      RECT 477.500000 0.000000 478.970000 0.630000 ;
      RECT 475.605000 0.000000 477.080000 0.630000 ;
      RECT 473.710000 0.000000 475.185000 0.630000 ;
      RECT 471.815000 0.000000 473.290000 0.630000 ;
      RECT 469.920000 0.000000 471.395000 0.630000 ;
      RECT 468.030000 0.000000 469.500000 0.630000 ;
      RECT 466.135000 0.000000 467.610000 0.630000 ;
      RECT 464.240000 0.000000 465.715000 0.630000 ;
      RECT 462.345000 0.000000 463.820000 0.630000 ;
      RECT 460.450000 0.000000 461.925000 0.630000 ;
      RECT 458.560000 0.000000 460.030000 0.630000 ;
      RECT 456.665000 0.000000 458.140000 0.630000 ;
      RECT 454.770000 0.000000 456.245000 0.630000 ;
      RECT 452.875000 0.000000 454.350000 0.630000 ;
      RECT 450.980000 0.000000 452.455000 0.630000 ;
      RECT 449.090000 0.000000 450.560000 0.630000 ;
      RECT 447.195000 0.000000 448.670000 0.630000 ;
      RECT 445.300000 0.000000 446.775000 0.630000 ;
      RECT 443.405000 0.000000 444.880000 0.630000 ;
      RECT 441.510000 0.000000 442.985000 0.630000 ;
      RECT 439.620000 0.000000 441.090000 0.630000 ;
      RECT 437.725000 0.000000 439.200000 0.630000 ;
      RECT 435.830000 0.000000 437.305000 0.630000 ;
      RECT 433.935000 0.000000 435.410000 0.630000 ;
      RECT 432.040000 0.000000 433.515000 0.630000 ;
      RECT 430.150000 0.000000 431.620000 0.630000 ;
      RECT 428.255000 0.000000 429.730000 0.630000 ;
      RECT 426.360000 0.000000 427.835000 0.630000 ;
      RECT 424.465000 0.000000 425.940000 0.630000 ;
      RECT 422.570000 0.000000 424.045000 0.630000 ;
      RECT 420.680000 0.000000 422.150000 0.630000 ;
      RECT 418.785000 0.000000 420.260000 0.630000 ;
      RECT 416.890000 0.000000 418.365000 0.630000 ;
      RECT 414.995000 0.000000 416.470000 0.630000 ;
      RECT 413.100000 0.000000 414.575000 0.630000 ;
      RECT 411.210000 0.000000 412.680000 0.630000 ;
      RECT 409.315000 0.000000 410.790000 0.630000 ;
      RECT 407.420000 0.000000 408.895000 0.630000 ;
      RECT 405.525000 0.000000 407.000000 0.630000 ;
      RECT 403.630000 0.000000 405.105000 0.630000 ;
      RECT 401.740000 0.000000 403.210000 0.630000 ;
      RECT 399.845000 0.000000 401.320000 0.630000 ;
      RECT 397.950000 0.000000 399.425000 0.630000 ;
      RECT 396.055000 0.000000 397.530000 0.630000 ;
      RECT 394.160000 0.000000 395.635000 0.630000 ;
      RECT 392.270000 0.000000 393.740000 0.630000 ;
      RECT 390.375000 0.000000 391.850000 0.630000 ;
      RECT 388.480000 0.000000 389.955000 0.630000 ;
      RECT 386.585000 0.000000 388.060000 0.630000 ;
      RECT 384.690000 0.000000 386.165000 0.630000 ;
      RECT 382.800000 0.000000 384.270000 0.630000 ;
      RECT 380.905000 0.000000 382.380000 0.630000 ;
      RECT 379.010000 0.000000 380.485000 0.630000 ;
      RECT 377.115000 0.000000 378.590000 0.630000 ;
      RECT 375.220000 0.000000 376.695000 0.630000 ;
      RECT 373.330000 0.000000 374.800000 0.630000 ;
      RECT 371.435000 0.000000 372.910000 0.630000 ;
      RECT 369.540000 0.000000 371.015000 0.630000 ;
      RECT 367.645000 0.000000 369.120000 0.630000 ;
      RECT 365.750000 0.000000 367.225000 0.630000 ;
      RECT 363.860000 0.000000 365.330000 0.630000 ;
      RECT 361.965000 0.000000 363.440000 0.630000 ;
      RECT 360.070000 0.000000 361.545000 0.630000 ;
      RECT 358.175000 0.000000 359.650000 0.630000 ;
      RECT 356.280000 0.000000 357.755000 0.630000 ;
      RECT 354.390000 0.000000 355.860000 0.630000 ;
      RECT 352.495000 0.000000 353.970000 0.630000 ;
      RECT 350.600000 0.000000 352.075000 0.630000 ;
      RECT 348.705000 0.000000 350.180000 0.630000 ;
      RECT 346.810000 0.000000 348.285000 0.630000 ;
      RECT 344.920000 0.000000 346.390000 0.630000 ;
      RECT 343.025000 0.000000 344.500000 0.630000 ;
      RECT 341.130000 0.000000 342.605000 0.630000 ;
      RECT 339.235000 0.000000 340.710000 0.630000 ;
      RECT 337.340000 0.000000 338.815000 0.630000 ;
      RECT 335.450000 0.000000 336.920000 0.630000 ;
      RECT 333.555000 0.000000 335.030000 0.630000 ;
      RECT 331.660000 0.000000 333.135000 0.630000 ;
      RECT 329.765000 0.000000 331.240000 0.630000 ;
      RECT 327.870000 0.000000 329.345000 0.630000 ;
      RECT 325.980000 0.000000 327.450000 0.630000 ;
      RECT 324.085000 0.000000 325.560000 0.630000 ;
      RECT 322.190000 0.000000 323.665000 0.630000 ;
      RECT 320.295000 0.000000 321.770000 0.630000 ;
      RECT 318.400000 0.000000 319.875000 0.630000 ;
      RECT 316.510000 0.000000 317.980000 0.630000 ;
      RECT 314.615000 0.000000 316.090000 0.630000 ;
      RECT 312.720000 0.000000 314.195000 0.630000 ;
      RECT 310.825000 0.000000 312.300000 0.630000 ;
      RECT 308.930000 0.000000 310.405000 0.630000 ;
      RECT 307.040000 0.000000 308.510000 0.630000 ;
      RECT 305.145000 0.000000 306.620000 0.630000 ;
      RECT 303.250000 0.000000 304.725000 0.630000 ;
      RECT 301.355000 0.000000 302.830000 0.630000 ;
      RECT 299.460000 0.000000 300.935000 0.630000 ;
      RECT 297.570000 0.000000 299.040000 0.630000 ;
      RECT 295.675000 0.000000 297.150000 0.630000 ;
      RECT 293.780000 0.000000 295.255000 0.630000 ;
      RECT 291.885000 0.000000 293.360000 0.630000 ;
      RECT 289.990000 0.000000 291.465000 0.630000 ;
      RECT 288.100000 0.000000 289.570000 0.630000 ;
      RECT 286.205000 0.000000 287.680000 0.630000 ;
      RECT 284.310000 0.000000 285.785000 0.630000 ;
      RECT 282.415000 0.000000 283.890000 0.630000 ;
      RECT 280.520000 0.000000 281.995000 0.630000 ;
      RECT 278.630000 0.000000 280.100000 0.630000 ;
      RECT 276.735000 0.000000 278.210000 0.630000 ;
      RECT 274.840000 0.000000 276.315000 0.630000 ;
      RECT 272.945000 0.000000 274.420000 0.630000 ;
      RECT 271.050000 0.000000 272.525000 0.630000 ;
      RECT 269.160000 0.000000 270.630000 0.630000 ;
      RECT 267.265000 0.000000 268.740000 0.630000 ;
      RECT 265.370000 0.000000 266.845000 0.630000 ;
      RECT 263.475000 0.000000 264.950000 0.630000 ;
      RECT 261.580000 0.000000 263.055000 0.630000 ;
      RECT 259.690000 0.000000 261.160000 0.630000 ;
      RECT 257.795000 0.000000 259.270000 0.630000 ;
      RECT 255.900000 0.000000 257.375000 0.630000 ;
      RECT 254.005000 0.000000 255.480000 0.630000 ;
      RECT 252.110000 0.000000 253.585000 0.630000 ;
      RECT 250.220000 0.000000 251.690000 0.630000 ;
      RECT 248.325000 0.000000 249.800000 0.630000 ;
      RECT 246.430000 0.000000 247.905000 0.630000 ;
      RECT 244.535000 0.000000 246.010000 0.630000 ;
      RECT 242.640000 0.000000 244.115000 0.630000 ;
      RECT 240.750000 0.000000 242.220000 0.630000 ;
      RECT 238.855000 0.000000 240.330000 0.630000 ;
      RECT 236.960000 0.000000 238.435000 0.630000 ;
      RECT 235.065000 0.000000 236.540000 0.630000 ;
      RECT 233.170000 0.000000 234.645000 0.630000 ;
      RECT 231.280000 0.000000 232.750000 0.630000 ;
      RECT 229.385000 0.000000 230.860000 0.630000 ;
      RECT 227.490000 0.000000 228.965000 0.630000 ;
      RECT 225.595000 0.000000 227.070000 0.630000 ;
      RECT 223.700000 0.000000 225.175000 0.630000 ;
      RECT 221.810000 0.000000 223.280000 0.630000 ;
      RECT 219.915000 0.000000 221.390000 0.630000 ;
      RECT 218.020000 0.000000 219.495000 0.630000 ;
      RECT 216.125000 0.000000 217.600000 0.630000 ;
      RECT 214.230000 0.000000 215.705000 0.630000 ;
      RECT 212.340000 0.000000 213.810000 0.630000 ;
      RECT 210.445000 0.000000 211.920000 0.630000 ;
      RECT 208.550000 0.000000 210.025000 0.630000 ;
      RECT 206.655000 0.000000 208.130000 0.630000 ;
      RECT 204.760000 0.000000 206.235000 0.630000 ;
      RECT 202.870000 0.000000 204.340000 0.630000 ;
      RECT 200.975000 0.000000 202.450000 0.630000 ;
      RECT 199.080000 0.000000 200.555000 0.630000 ;
      RECT 197.185000 0.000000 198.660000 0.630000 ;
      RECT 195.290000 0.000000 196.765000 0.630000 ;
      RECT 193.400000 0.000000 194.870000 0.630000 ;
      RECT 191.505000 0.000000 192.980000 0.630000 ;
      RECT 189.610000 0.000000 191.085000 0.630000 ;
      RECT 187.715000 0.000000 189.190000 0.630000 ;
      RECT 185.820000 0.000000 187.295000 0.630000 ;
      RECT 183.930000 0.000000 185.400000 0.630000 ;
      RECT 182.035000 0.000000 183.510000 0.630000 ;
      RECT 180.140000 0.000000 181.615000 0.630000 ;
      RECT 178.245000 0.000000 179.720000 0.630000 ;
      RECT 176.350000 0.000000 177.825000 0.630000 ;
      RECT 174.460000 0.000000 175.930000 0.630000 ;
      RECT 172.565000 0.000000 174.040000 0.630000 ;
      RECT 170.670000 0.000000 172.145000 0.630000 ;
      RECT 168.775000 0.000000 170.250000 0.630000 ;
      RECT 166.880000 0.000000 168.355000 0.630000 ;
      RECT 164.990000 0.000000 166.460000 0.630000 ;
      RECT 163.095000 0.000000 164.570000 0.630000 ;
      RECT 161.200000 0.000000 162.675000 0.630000 ;
      RECT 159.305000 0.000000 160.780000 0.630000 ;
      RECT 157.410000 0.000000 158.885000 0.630000 ;
      RECT 155.520000 0.000000 156.990000 0.630000 ;
      RECT 153.625000 0.000000 155.100000 0.630000 ;
      RECT 151.730000 0.000000 153.205000 0.630000 ;
      RECT 149.835000 0.000000 151.310000 0.630000 ;
      RECT 147.940000 0.000000 149.415000 0.630000 ;
      RECT 146.050000 0.000000 147.520000 0.630000 ;
      RECT 144.155000 0.000000 145.630000 0.630000 ;
      RECT 142.260000 0.000000 143.735000 0.630000 ;
      RECT 140.365000 0.000000 141.840000 0.630000 ;
      RECT 138.470000 0.000000 139.945000 0.630000 ;
      RECT 136.580000 0.000000 138.050000 0.630000 ;
      RECT 134.685000 0.000000 136.160000 0.630000 ;
      RECT 132.790000 0.000000 134.265000 0.630000 ;
      RECT 130.895000 0.000000 132.370000 0.630000 ;
      RECT 129.000000 0.000000 130.475000 0.630000 ;
      RECT 127.110000 0.000000 128.580000 0.630000 ;
      RECT 125.215000 0.000000 126.690000 0.630000 ;
      RECT 123.320000 0.000000 124.795000 0.630000 ;
      RECT 121.425000 0.000000 122.900000 0.630000 ;
      RECT 119.530000 0.000000 121.005000 0.630000 ;
      RECT 117.640000 0.000000 119.110000 0.630000 ;
      RECT 115.745000 0.000000 117.220000 0.630000 ;
      RECT 113.850000 0.000000 115.325000 0.630000 ;
      RECT 111.955000 0.000000 113.430000 0.630000 ;
      RECT 110.060000 0.000000 111.535000 0.630000 ;
      RECT 108.170000 0.000000 109.640000 0.630000 ;
      RECT 106.275000 0.000000 107.750000 0.630000 ;
      RECT 104.380000 0.000000 105.855000 0.630000 ;
      RECT 102.485000 0.000000 103.960000 0.630000 ;
      RECT 100.590000 0.000000 102.065000 0.630000 ;
      RECT 98.700000 0.000000 100.170000 0.630000 ;
      RECT 96.805000 0.000000 98.280000 0.630000 ;
      RECT 94.910000 0.000000 96.385000 0.630000 ;
      RECT 93.015000 0.000000 94.490000 0.630000 ;
      RECT 91.120000 0.000000 92.595000 0.630000 ;
      RECT 89.230000 0.000000 90.700000 0.630000 ;
      RECT 87.335000 0.000000 88.810000 0.630000 ;
      RECT 85.440000 0.000000 86.915000 0.630000 ;
      RECT 83.545000 0.000000 85.020000 0.630000 ;
      RECT 81.650000 0.000000 83.125000 0.630000 ;
      RECT 79.760000 0.000000 81.230000 0.630000 ;
      RECT 77.865000 0.000000 79.340000 0.630000 ;
      RECT 75.970000 0.000000 77.445000 0.630000 ;
      RECT 74.075000 0.000000 75.550000 0.630000 ;
      RECT 72.180000 0.000000 73.655000 0.630000 ;
      RECT 70.290000 0.000000 71.760000 0.630000 ;
      RECT 68.395000 0.000000 69.870000 0.630000 ;
      RECT 66.500000 0.000000 67.975000 0.630000 ;
      RECT 64.605000 0.000000 66.080000 0.630000 ;
      RECT 62.710000 0.000000 64.185000 0.630000 ;
      RECT 60.820000 0.000000 62.290000 0.630000 ;
      RECT 58.925000 0.000000 60.400000 0.630000 ;
      RECT 57.030000 0.000000 58.505000 0.630000 ;
      RECT 55.135000 0.000000 56.610000 0.630000 ;
      RECT 53.240000 0.000000 54.715000 0.630000 ;
      RECT 51.350000 0.000000 52.820000 0.630000 ;
      RECT 49.455000 0.000000 50.930000 0.630000 ;
      RECT 47.560000 0.000000 49.035000 0.630000 ;
      RECT 45.665000 0.000000 47.140000 0.630000 ;
      RECT 43.770000 0.000000 45.245000 0.630000 ;
      RECT 41.880000 0.000000 43.350000 0.630000 ;
      RECT 39.985000 0.000000 41.460000 0.630000 ;
      RECT 38.090000 0.000000 39.565000 0.630000 ;
      RECT 36.195000 0.000000 37.670000 0.630000 ;
      RECT 34.300000 0.000000 35.775000 0.630000 ;
      RECT 32.410000 0.000000 33.880000 0.630000 ;
      RECT 30.515000 0.000000 31.990000 0.630000 ;
      RECT 28.620000 0.000000 30.095000 0.630000 ;
      RECT 26.725000 0.000000 28.200000 0.630000 ;
      RECT 24.830000 0.000000 26.305000 0.630000 ;
      RECT 22.940000 0.000000 24.410000 0.630000 ;
      RECT 21.045000 0.000000 22.520000 0.630000 ;
      RECT 19.150000 0.000000 20.625000 0.630000 ;
      RECT 17.255000 0.000000 18.730000 0.630000 ;
      RECT 15.360000 0.000000 16.835000 0.630000 ;
      RECT 13.470000 0.000000 14.940000 0.630000 ;
      RECT 11.575000 0.000000 13.050000 0.630000 ;
      RECT 9.680000 0.000000 11.155000 0.630000 ;
      RECT 7.785000 0.000000 9.260000 0.630000 ;
      RECT 5.890000 0.000000 7.365000 0.630000 ;
      RECT 4.000000 0.000000 5.470000 0.630000 ;
      RECT 2.105000 0.000000 3.580000 0.630000 ;
      RECT 1.360000 0.000000 1.685000 0.630000 ;
      RECT 0.000000 0.000000 0.940000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 920.330000 926.440000 923.440000 ;
      RECT 1.100000 919.430000 925.340000 920.330000 ;
      RECT 0.000000 902.890000 926.440000 919.430000 ;
      RECT 0.000000 901.990000 925.340000 902.890000 ;
      RECT 0.000000 901.330000 926.440000 901.990000 ;
      RECT 1.100000 900.430000 926.440000 901.330000 ;
      RECT 0.000000 881.905000 926.440000 900.430000 ;
      RECT 0.000000 881.005000 925.340000 881.905000 ;
      RECT 0.000000 878.810000 926.440000 881.005000 ;
      RECT 1.100000 877.910000 926.440000 878.810000 ;
      RECT 0.000000 860.915000 926.440000 877.910000 ;
      RECT 0.000000 860.015000 925.340000 860.915000 ;
      RECT 0.000000 856.285000 926.440000 860.015000 ;
      RECT 1.100000 855.385000 926.440000 856.285000 ;
      RECT 0.000000 839.930000 926.440000 855.385000 ;
      RECT 0.000000 839.030000 925.340000 839.930000 ;
      RECT 0.000000 833.765000 926.440000 839.030000 ;
      RECT 1.100000 832.865000 926.440000 833.765000 ;
      RECT 0.000000 818.945000 926.440000 832.865000 ;
      RECT 0.000000 818.045000 925.340000 818.945000 ;
      RECT 0.000000 811.240000 926.440000 818.045000 ;
      RECT 1.100000 810.340000 926.440000 811.240000 ;
      RECT 0.000000 797.955000 926.440000 810.340000 ;
      RECT 0.000000 797.055000 925.340000 797.955000 ;
      RECT 0.000000 788.720000 926.440000 797.055000 ;
      RECT 1.100000 787.820000 926.440000 788.720000 ;
      RECT 0.000000 776.970000 926.440000 787.820000 ;
      RECT 0.000000 776.070000 925.340000 776.970000 ;
      RECT 0.000000 766.200000 926.440000 776.070000 ;
      RECT 1.100000 765.300000 926.440000 766.200000 ;
      RECT 0.000000 755.980000 926.440000 765.300000 ;
      RECT 0.000000 755.080000 925.340000 755.980000 ;
      RECT 0.000000 743.675000 926.440000 755.080000 ;
      RECT 1.100000 742.775000 926.440000 743.675000 ;
      RECT 0.000000 734.995000 926.440000 742.775000 ;
      RECT 0.000000 734.095000 925.340000 734.995000 ;
      RECT 0.000000 721.155000 926.440000 734.095000 ;
      RECT 1.100000 720.255000 926.440000 721.155000 ;
      RECT 0.000000 714.010000 926.440000 720.255000 ;
      RECT 0.000000 713.110000 925.340000 714.010000 ;
      RECT 0.000000 698.630000 926.440000 713.110000 ;
      RECT 1.100000 697.730000 926.440000 698.630000 ;
      RECT 0.000000 693.020000 926.440000 697.730000 ;
      RECT 0.000000 692.120000 925.340000 693.020000 ;
      RECT 0.000000 676.110000 926.440000 692.120000 ;
      RECT 1.100000 675.210000 926.440000 676.110000 ;
      RECT 0.000000 672.035000 926.440000 675.210000 ;
      RECT 0.000000 671.135000 925.340000 672.035000 ;
      RECT 0.000000 653.590000 926.440000 671.135000 ;
      RECT 1.100000 652.690000 926.440000 653.590000 ;
      RECT 0.000000 651.045000 926.440000 652.690000 ;
      RECT 0.000000 650.145000 925.340000 651.045000 ;
      RECT 0.000000 631.065000 926.440000 650.145000 ;
      RECT 1.100000 630.165000 926.440000 631.065000 ;
      RECT 0.000000 630.060000 926.440000 630.165000 ;
      RECT 0.000000 629.160000 925.340000 630.060000 ;
      RECT 0.000000 609.075000 926.440000 629.160000 ;
      RECT 0.000000 608.545000 925.340000 609.075000 ;
      RECT 1.100000 608.175000 925.340000 608.545000 ;
      RECT 1.100000 607.645000 926.440000 608.175000 ;
      RECT 0.000000 588.085000 926.440000 607.645000 ;
      RECT 0.000000 587.185000 925.340000 588.085000 ;
      RECT 0.000000 586.020000 926.440000 587.185000 ;
      RECT 1.100000 585.120000 926.440000 586.020000 ;
      RECT 0.000000 567.100000 926.440000 585.120000 ;
      RECT 0.000000 566.200000 925.340000 567.100000 ;
      RECT 0.000000 563.500000 926.440000 566.200000 ;
      RECT 1.100000 562.600000 926.440000 563.500000 ;
      RECT 0.000000 546.110000 926.440000 562.600000 ;
      RECT 0.000000 545.210000 925.340000 546.110000 ;
      RECT 0.000000 540.980000 926.440000 545.210000 ;
      RECT 1.100000 540.080000 926.440000 540.980000 ;
      RECT 0.000000 525.125000 926.440000 540.080000 ;
      RECT 0.000000 524.225000 925.340000 525.125000 ;
      RECT 0.000000 518.455000 926.440000 524.225000 ;
      RECT 1.100000 517.555000 926.440000 518.455000 ;
      RECT 0.000000 504.140000 926.440000 517.555000 ;
      RECT 0.000000 503.240000 925.340000 504.140000 ;
      RECT 0.000000 495.935000 926.440000 503.240000 ;
      RECT 1.100000 495.035000 926.440000 495.935000 ;
      RECT 0.000000 483.150000 926.440000 495.035000 ;
      RECT 0.000000 482.250000 925.340000 483.150000 ;
      RECT 0.000000 473.410000 926.440000 482.250000 ;
      RECT 1.100000 472.510000 926.440000 473.410000 ;
      RECT 0.000000 462.165000 926.440000 472.510000 ;
      RECT 0.000000 461.265000 925.340000 462.165000 ;
      RECT 0.000000 450.890000 926.440000 461.265000 ;
      RECT 1.100000 449.990000 926.440000 450.890000 ;
      RECT 0.000000 441.175000 926.440000 449.990000 ;
      RECT 0.000000 440.275000 925.340000 441.175000 ;
      RECT 0.000000 428.370000 926.440000 440.275000 ;
      RECT 1.100000 427.470000 926.440000 428.370000 ;
      RECT 0.000000 420.190000 926.440000 427.470000 ;
      RECT 0.000000 419.290000 925.340000 420.190000 ;
      RECT 0.000000 405.845000 926.440000 419.290000 ;
      RECT 1.100000 404.945000 926.440000 405.845000 ;
      RECT 0.000000 399.205000 926.440000 404.945000 ;
      RECT 0.000000 398.305000 925.340000 399.205000 ;
      RECT 0.000000 383.325000 926.440000 398.305000 ;
      RECT 1.100000 382.425000 926.440000 383.325000 ;
      RECT 0.000000 378.215000 926.440000 382.425000 ;
      RECT 0.000000 377.315000 925.340000 378.215000 ;
      RECT 0.000000 360.800000 926.440000 377.315000 ;
      RECT 1.100000 359.900000 926.440000 360.800000 ;
      RECT 0.000000 357.230000 926.440000 359.900000 ;
      RECT 0.000000 356.330000 925.340000 357.230000 ;
      RECT 0.000000 338.280000 926.440000 356.330000 ;
      RECT 1.100000 337.380000 926.440000 338.280000 ;
      RECT 0.000000 336.240000 926.440000 337.380000 ;
      RECT 0.000000 335.340000 925.340000 336.240000 ;
      RECT 0.000000 315.760000 926.440000 335.340000 ;
      RECT 1.100000 315.255000 926.440000 315.760000 ;
      RECT 1.100000 314.860000 925.340000 315.255000 ;
      RECT 0.000000 314.355000 925.340000 314.860000 ;
      RECT 0.000000 294.270000 926.440000 314.355000 ;
      RECT 0.000000 293.370000 925.340000 294.270000 ;
      RECT 0.000000 293.235000 926.440000 293.370000 ;
      RECT 1.100000 292.335000 926.440000 293.235000 ;
      RECT 0.000000 273.280000 926.440000 292.335000 ;
      RECT 0.000000 272.380000 925.340000 273.280000 ;
      RECT 0.000000 270.715000 926.440000 272.380000 ;
      RECT 1.100000 269.815000 926.440000 270.715000 ;
      RECT 0.000000 252.295000 926.440000 269.815000 ;
      RECT 0.000000 251.395000 925.340000 252.295000 ;
      RECT 0.000000 248.190000 926.440000 251.395000 ;
      RECT 1.100000 247.290000 926.440000 248.190000 ;
      RECT 0.000000 231.305000 926.440000 247.290000 ;
      RECT 0.000000 230.405000 925.340000 231.305000 ;
      RECT 0.000000 225.670000 926.440000 230.405000 ;
      RECT 1.100000 224.770000 926.440000 225.670000 ;
      RECT 0.000000 210.320000 926.440000 224.770000 ;
      RECT 0.000000 209.420000 925.340000 210.320000 ;
      RECT 0.000000 203.150000 926.440000 209.420000 ;
      RECT 1.100000 202.250000 926.440000 203.150000 ;
      RECT 0.000000 189.335000 926.440000 202.250000 ;
      RECT 0.000000 188.435000 925.340000 189.335000 ;
      RECT 0.000000 180.625000 926.440000 188.435000 ;
      RECT 1.100000 179.725000 926.440000 180.625000 ;
      RECT 0.000000 168.345000 926.440000 179.725000 ;
      RECT 0.000000 167.445000 925.340000 168.345000 ;
      RECT 0.000000 158.105000 926.440000 167.445000 ;
      RECT 1.100000 157.205000 926.440000 158.105000 ;
      RECT 0.000000 147.360000 926.440000 157.205000 ;
      RECT 0.000000 146.460000 925.340000 147.360000 ;
      RECT 0.000000 135.580000 926.440000 146.460000 ;
      RECT 1.100000 134.680000 926.440000 135.580000 ;
      RECT 0.000000 126.370000 926.440000 134.680000 ;
      RECT 0.000000 125.470000 925.340000 126.370000 ;
      RECT 0.000000 113.060000 926.440000 125.470000 ;
      RECT 1.100000 112.160000 926.440000 113.060000 ;
      RECT 0.000000 105.385000 926.440000 112.160000 ;
      RECT 0.000000 104.485000 925.340000 105.385000 ;
      RECT 0.000000 90.540000 926.440000 104.485000 ;
      RECT 1.100000 89.640000 926.440000 90.540000 ;
      RECT 0.000000 84.400000 926.440000 89.640000 ;
      RECT 0.000000 83.500000 925.340000 84.400000 ;
      RECT 0.000000 68.015000 926.440000 83.500000 ;
      RECT 1.100000 67.115000 926.440000 68.015000 ;
      RECT 0.000000 63.410000 926.440000 67.115000 ;
      RECT 0.000000 62.510000 925.340000 63.410000 ;
      RECT 0.000000 45.495000 926.440000 62.510000 ;
      RECT 1.100000 44.595000 926.440000 45.495000 ;
      RECT 0.000000 42.425000 926.440000 44.595000 ;
      RECT 0.000000 41.525000 925.340000 42.425000 ;
      RECT 0.000000 22.970000 926.440000 41.525000 ;
      RECT 1.100000 22.070000 926.440000 22.970000 ;
      RECT 0.000000 21.435000 926.440000 22.070000 ;
      RECT 0.000000 20.535000 925.340000 21.435000 ;
      RECT 0.000000 15.700000 926.440000 20.535000 ;
      RECT 1.100000 14.800000 926.440000 15.700000 ;
      RECT 0.000000 10.820000 926.440000 14.800000 ;
      RECT 1.100000 9.920000 926.440000 10.820000 ;
      RECT 0.000000 5.940000 926.440000 9.920000 ;
      RECT 1.100000 5.330000 926.440000 5.940000 ;
      RECT 1.100000 5.040000 925.340000 5.330000 ;
      RECT 0.000000 4.430000 925.340000 5.040000 ;
      RECT 0.000000 1.100000 926.440000 4.430000 ;
      RECT 1.140000 0.000000 926.440000 1.100000 ;
      RECT 0.000000 0.000000 0.240000 1.100000 ;
    LAYER met4 ;
      RECT 0.000000 921.640000 926.440000 923.440000 ;
      RECT 4.360000 917.640000 922.080000 921.640000 ;
      RECT 920.680000 5.800000 922.080000 917.640000 ;
      RECT 8.360000 5.800000 918.080000 917.640000 ;
      RECT 4.360000 5.800000 5.760000 917.640000 ;
      RECT 924.680000 1.800000 926.440000 921.640000 ;
      RECT 4.360000 1.800000 922.080000 5.800000 ;
      RECT 0.000000 1.800000 1.760000 921.640000 ;
      RECT 0.000000 0.000000 926.440000 1.800000 ;
  END
END user_proj_example

END LIBRARY
